/*=============================================================================
// RUIJIE IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS"
// SOLELY FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR
// RUIJIE DEVICES.  BY PROVIDING THIS DESIGN, CODE, OR INFORMATION
// AS ONE POSSIBLE IMPLEMENTATION OF THIS FEATURE, APPLICATION
// OR STANDARD, RUIJIE IS MAKING NO REPRESENTATION THAT THIS
// IMPLEMENTATION IS FREE FROM ANY CLAIMS OF INFRINGEMENT,
// AND YOU ARE RESPONSIBLE FOR OBTAINING ANY RIGHTS YOU MAY REQUIRE
// FOR YOUR IMPLEMENTATION.  RUIJIE EXPRESSLY DISCLAIMS ANY
// WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE
// IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR
// REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF
// INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS
// FOR A PARTICULAR PURPOSE.
// (c) Copyright 2007 RUIJIE, Inc.
// All rights reserved.

//============================================================================
//     FileName: pcie_tlp_monitor.sv
//         Desc:  
//       Author: lixu
//        Email: lixu@ruijie.com.cn
//     HomePage: http://www.ruijie.com.cn
//      Version: 0.0.1
//   LastChange: 2016-04-21 17:47:06
//      History:
//============================================================================*/
`ifndef PCIE_TLP_MONITOR__SV
`define PCIE_TLP_MONITOR__SV

class pcie_tlp_monitor extends uvm_monitor;
  
	`SET_CLASSID
	pcie_tlp_cfg  m_cfg;
	abstract_if m_pcie_tlp_vif;
	uvm_analysis_port     #(pcie_tlp_pkt)  mon_analysis_port; 
	uvm_analysis_export   #(pcie_tlp_pkt)  drv2mon_export; 
	uvm_tlm_analysis_fifo #(pcie_tlp_pkt)  drv2mon_afifo;
	pcie_tlp_pkt drv2mon_req_aq[int][$];
	
	uvm_thread reset_handler;
	local uvm_thread_imp#(pcie_tlp_monitor) reset_export;

	`uvm_component_utils_begin(pcie_tlp_monitor)
        `uvm_field_object(reset_handler, UVM_DEFAULT|UVM_REFERENCE)
	`uvm_component_utils_end

	function new (string name = "pcie_tlp_monitor", uvm_component parent = null);
		super.new(name, parent);
		reset_export = new("reset_export", this);
		mon_analysis_port = new("mon_analysis_port", this);
		drv2mon_export = new("mon_export", this);
		drv2mon_afifo = new("drv2mon_afifo", this);
	endfunction: new

	extern virtual function void build_phase(uvm_phase phase);
	extern virtual function void connect_phase(uvm_phase phase);
	extern virtual task main_phase(uvm_phase phase);
	extern virtual task clean_up();
    extern virtual task main_phase_new(uvm_phase phase);
	extern virtual task collect_transactions();

endclass: pcie_tlp_monitor

function void pcie_tlp_monitor::build_phase(input uvm_phase phase);
	super.build_phase(phase);
	if (!uvm_config_db#(pcie_tlp_cfg)::get(this, "", "pcie_tlp_cfg", m_cfg)) begin
		`uvm_fatal(CLASSID, "Failed to Grab pcie_tlp_cfg from Config DB")
	end
	if (!uvm_config_db#(abstract_if)::get(this, "", "PCIE_TLP_IF", m_pcie_tlp_vif)) begin
		`uvm_fatal(CLASSID, "Failed to Grab pcie_tlp_if from Config DB")
	end

	if (reset_handler == null) begin 
		if (!uvm_config_db#(uvm_thread)::get(this, "", "reset_handler", reset_handler))
			`uvm_fatal(CLASSID, "reset_handler must be specified")
	end
	reset_handler.register(reset_export, uvm_thread_pkg::default_map);
endfunction: build_phase


function void pcie_tlp_monitor::connect_phase(input uvm_phase phase);
	drv2mon_export.connect(drv2mon_afifo.analysis_export); 
endfunction: connect_phase

task pcie_tlp_monitor::main_phase(uvm_phase phase);
endtask: main_phase

task pcie_tlp_monitor::clean_up();
	`uvm_info(CLASSID, "CLEANING...........................", UVM_MEDIUM)
	disable collect_transactions;
	m_pcie_tlp_vif.clean_up();
endtask : clean_up

task pcie_tlp_monitor::main_phase_new(uvm_phase phase);
	`uvm_info(CLASSID, "Now Collecting Transactions.....................", UVM_MEDIUM)
	fork
		forever begin 
		    pcie_tlp_pkt req;
		    drv2mon_afifo.get(req);
			if(req.pcie_tlp_type == MRD) begin 
				drv2mon_req_aq[{req.req_id,req.tag}].push_back(req);
			end
			else if(req.pcie_tlp_type inside {MRDLK,IORD,IOWR,CFGRD0,CFGRD1,CFGWR0,CFGWR1}) begin 
				`uvm_fatal(CLASSID,$sformatf("Can not support TLP TYPE[%p]!",req.pcie_tlp_type))
			end
		end
	    collect_transactions();
    join
endtask : main_phase_new

task pcie_tlp_monitor::collect_transactions();
	uvm_sequence_item mon_item;
	pcie_tlp_pkt m_pkt;
	bit [7:0] data_q[int][$];
	bit finish[int] = '{default:0};
	int pid;
    forever begin 
		m_pcie_tlp_vif.recvPkt(mon_item);
		$cast(m_pkt,mon_item.clone());
		//#################################################################
		m_pkt.fmt = m_pkt.pcie_tlp_data[0][6:5];
		m_pkt.typ = m_pkt.pcie_tlp_data[0][4:0];
		if(m_pkt.fmt == 2'b10 && m_pkt.typ == 5'b01010) begin 
			m_pkt.pcie_tlp_type = CPLD;
			m_pkt.is_cpl_op = 1;
			m_pkt.is_with_data = 1;
		end
		else
			`uvm_fatal(CLASSID,$sformatf("You recvPkt has wrong type: ----->\n%0s",m_pkt.sprint()))
		m_pkt.tc = m_pkt.pcie_tlp_data[1][6:4];
		m_pkt.td = m_pkt.pcie_tlp_data[2][7];
		m_pkt.ep = m_pkt.pcie_tlp_data[2][6];
		m_pkt.attr = m_pkt.pcie_tlp_data[2][5:4];
		m_pkt.length = {m_pkt.pcie_tlp_data[2][1:0],m_pkt.pcie_tlp_data[3]};
		m_pkt.cpl_id = {m_pkt.pcie_tlp_data[4],m_pkt.pcie_tlp_data[5]};
		m_pkt.cpl_st = m_pkt.pcie_tlp_data[6][7:5];
		m_pkt.bcm = m_pkt.pcie_tlp_data[6][4];
		m_pkt.byte_cnt = {m_pkt.pcie_tlp_data[6][3:0],m_pkt.pcie_tlp_data[7]};
		m_pkt.req_id = {m_pkt.pcie_tlp_data[8],m_pkt.pcie_tlp_data[9]};
		m_pkt.tag = m_pkt.pcie_tlp_data[10];
		m_pkt.lower_addr = m_pkt.pcie_tlp_data[11][6:0];
		m_pkt.pcie_tlp_data = m_pkt.pcie_tlp_data[12:$];
		pid = {m_pkt.req_id,m_pkt.tag};
		//#################################################################
		if(m_pkt.bcm == 1) 
			`uvm_fatal(CLASSID,$sformatf("You recvPkt has BCM == 1 : ----->\n%0s",m_pkt.sprint()))
		if(m_pkt.ep == 1)
			`uvm_fatal(CLASSID,$sformatf("You recvPkt has EP == 1 : ----->\n%0s",m_pkt.sprint()))
		if(m_pkt.cpl_st != 3'b0)
			`uvm_fatal(CLASSID,$sformatf("You recvPkt has wrong cpl_st: ----->\n%0s",m_pkt.sprint()))
		if(m_pkt.pcie_tlp_data.size() == 0) begin 
			`uvm_fatal(CLASSID,$sformatf("You recvPkt has no payload: ----->\n%0s",m_pkt.sprint()))
		end
		else if(m_pkt.pcie_tlp_data.size()%4 != 0) begin 
			`uvm_fatal(CLASSID,$sformatf("You recvPkt payload not 1DW align!: ----->\n%0s",m_pkt.sprint()))
		end
		else if(m_pkt.pcie_tlp_data.size() != m_pkt.length*4 ) begin 
			`uvm_fatal(CLASSID,$sformatf("You recvPkt payload size != pcie tlp length!: ----->\n%0s",m_pkt.sprint()))
		end
		else if(m_pkt.pcie_tlp_data.size() > m_cfg.RCBLen)
			`uvm_fatal(CLASSID,$sformatf("You recvPkt payload size > RCB bytes(%0d): ----->\n%0s",m_cfg.RCBLen,m_pkt.sprint()))
		if(drv2mon_req_aq.exists(pid) == 0)
			`uvm_fatal(CLASSID,$sformatf("[%0p] You recvPkt has wrong req_id and tag[pid:%0d]: ----->\n%0s",drv2mon_req_aq,pid,m_pkt.sprint()))
		else begin 
			int m_len;
			int m_byte_cnt;
			m_len = (m_pkt.length == 0) ? 4096 : m_pkt.length*4;
			m_byte_cnt = (m_pkt.byte_cnt == 0) ? 4096 : m_pkt.byte_cnt;
			for(int i=0;i<m_pkt.lower_addr[1:0];i++)
				void'(m_pkt.pcie_tlp_data.pop_front());
			if(m_byte_cnt <= m_len - m_pkt.lower_addr[1:0]) begin  
				finish[pid] = 1;
				for(int i=0;i< (m_len-m_pkt.lower_addr[1:0]-m_byte_cnt);i++)
					void'(m_pkt.pcie_tlp_data.pop_back());
			end
			data_q[pid] = {data_q[pid],m_pkt.pcie_tlp_data};
			if(finish[pid] == 1) begin 
				m_pkt.up_payload = data_q[pid];
				`uvm_info(CLASSID,$sformatf("Collecting complete Transactions is:---->\n%0s",m_pkt.sprint()), UVM_LOW)
				mon_analysis_port.write(m_pkt);
				finish[pid] = 0;
				data_q[pid].delete();
				drv2mon_req_aq.delete(pid);
			end
		end
	end
endtask : collect_transactions


`endif 
