`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FCKIrZkL6ivqf5zjLHS3q/MkdL/7/0Z/hkXoQrTOSE7HwwZIvsnBFDcj/mBTegu27XTQxadKCSvK
x2ykjqRzAg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
YONXZlGJSwyjcPbDTGpOGB/2GtQF1uruwBEh2RVasgjmMFLP+tTDJosYv6focH2YUJahRcRXERUG
cJC0MlMi+kGTm0tk8Xv8WMGm6LMy02GziKe59R7emiZZsjD0LvzJqFeI6Z8h0UBtW8W5QD00oXV0
jNpUKPNqCN/M+m332wk=

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
vjhHVMisA6cYfenQOXi0SRkqAasXJO2lyhMl2nRNL43T173I2pZdXJDnqkswwSZL5SLnFIpo4sfJ
kXGzacxvyiVY+ZIZUPY57zDLaB8T28aREkWJC0ei4NanTF9T/kUmnvFQQKAILSQ5+01oJZ08psbA
FA6lYaa5Sijlp6FXpX4=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
GJikz3XiiG2RL5voVnIpuK9vfiQwZB20e18fB+zjU86CmTqP9Na517aYoUmVunuPN3SDhCcns804
dl5jQf+1vPHoe06XteeOnRk2K1YH2HTbGaPYNbbWffCJNX0L5sfwwe/9jZspP0fryN3EkgkAFL6V
OUrPVW1qj6rbUG4P53yMSDwGqBRhDfWODyiv5xLyoNGn9/84nu4JfbqB1OhnKvy2RKJUYQQP75Wq
3fig9BgUUU1CP/dFNy3KrST0OahdFtWyOcQ5OdobFFL8RdZdxR4Hfj7+vV7nnvXmdPD7sVVyKs30
LUlIv48CvY8UiR/4X0pGUJLGs9ri7SRChjLmjQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
V1X05JPVST6xVK1Gt2Rcuepz1Hs6GKbAcBGOvdq1Sgu1aFodQPWO1E/LyCQ5FugE6zt6UnociNdc
WGRbcMvIZMGXnpOEIWqOBYiKhGEuXXQwipKKyXYGCNyaAU7UyZlIp+FLR/68aBslfMuyIef0JNbF
lY0ZsXWaVWYbafvOLlhVCfB1Uid2PKOPP12YD8HP8PEwQJ21iDy7PYtTqYqrzL9kphpAyuEe700D
dKsWQaO8UlaKlLnF+Kf3xx8VRewN0CSys9+kwRsF33chqhOzzhncghNObvBD3jrrSAi0N81LcVrP
RtfiSTgGoWRPLT2s+FsurHl83m6k8mvQp79cUA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
us0vZr9iBhHgeLI5myrNrcGSg05Z2BOyMKL2HO1H/5Uwy3iXF25X6/cxkReNrDoKsXLBbs3c4+JH
1IVwFst40ZfUwubjHMjDrVutA2qfdfzx7jfGghaCMxYxejRqmCOoYyR63R2KNM0UfHJnFlRFVG46
obrgbB8KUiE7Intd0jZPgcPAc2UTrmo4VAklO2bUWyZxaR34m73Yren+QKhONAy8JRSqXMZyL1qk
zgQKwxm2xlVEGZOaOTHIRZ9peYZjDVPfGZPKzmn2gLrgu2bbEOlaNKxx0gARnKPI3Cx+YhLC6WrO
2BdLDiLrPCh/5Asgj94qkMb7O31gaYN4OY5T8A==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 135936)
`pragma protect data_block
ZgMYGaL+t7A4Ymtttu59itt0Ur/MeXFK62HhQRyKQk7F6w9CXVIdbFz4j8jyd6Dt6uxXKioU1gzw
gWH5XphDeLGQmVG+eh9sQfYKRATGq126L36g25sPailRUX9YivYCb4GgKexWdlr41fP8/1+c8s3P
v6KZ806HDt2DR5zsQjwXeGQ9WHzrnsq/l9OtIWDYaGEYOP/F/jkbVPXcj7MDdZKXIV+UsnDxc8Do
rS+1n7+sU3kuc6z9f/pbz89OVtXWdZxgOPbo/KFld9cDqcn+/RcMUe69qq0F+Wq2MYUVmosYN3SD
qg1PYj1wIQBmvtpxeSQDxZYI1bBiMt3ppJuMCF4HsPMZ6cO9D0h+t/mQTC5yisBd/PKmwv0vZnIk
rQyDXNdWbc5qSiFULIhFs1Iuk8Vz1RJDeeLqTiLh5jvPJ47Y/1FCjOsWKoseJ3vQ83K3HjyqPZMR
oSQTINoZYExawD7AGub3uaqQrEWoJEUDQWsfell+mPg/qt5LPRGmvS1/oOm40p+VTLDgKjqfjMf2
FO5v37pjX5fX7ciM3AcKwkfU2+4a6PrfEjSb9esKDsmPRn9pu55/EbYj2c2/WvxkdZhSfPaBmVlT
o9rGIANo3aNouAzN8LsQKvIN6rc5E/EBZ79kEOKwxLGBp4hDQnUKkYR1x9DVOdiwHFB/OZ4SA3cr
WQRblxoFNYPnEPmb5iG265+E+Ir/1omHwZ/S0n8Zoz+LNWbLtzjayismYUDbC6U/BraphmFJGbF8
QpcN+tgga3hql8w/LuTpFSW1o1H+W3sBkUDWDMzRy+qjUPhEW4c+abt/JuwFOeZTDwV98F9hHHLh
w5/At1/H1kN8N7YB8d/4LBx1yfhAQ9zsPAWJsbymUWjZ5Fy5xjtPO7Zlm1paUFk/WKcMyzYU2BVn
BWYZGT2DpdorJWS9w8r6AZpXIYV+jlX1bMGgXqds9LiC/aHWXMyx89PoZ8YDEI2oAL5l/6BQjlQ4
udKgYgtd9k1dQfVXQkdjo6/t8UOFyilc+0K1qmsbjctpAlYrLU5fjOxVstjgno8zcuR3XyFWb1dp
bIs075v9DSR3x5VuTfm4BcPHGTFe1eu4XCWkTOl1ounEgS2kpkazR6Os15iEMgNEzXTGXmrA6xwL
WmFH0BadxrjgPBDU5OM2jriw15zecNM0WiKtOn45uelHcewiHL/+7dPAI8QIIWkLHZCGqtY5Ttx6
ZzW/PKd0wfZiAtnIAUvqKtgTGBjngM/B5XwVFwkoy9k1dZ+XHa7bMJxdpt3fe73kPd8QTAraor8b
8iXKrChiZEB2a9IrrRUrn9v/cd1TPie/KvW1xPTsX8rXvDiiWkNOuYKhmyuoA3+Qgf2Cw0gNLux/
1/Fgz7UGJS3sCv9c7wmVUPJ/9eg2V9yx7x/aOUy8RXXOJebiT9+GfEArzTVWiAweT4+q2Z37YFPr
49fR9LScLqWpW8ARbcKUAMbUzgWyhMhyMsfWmQOV+zv4EmglYYb+zod2c5ST4SsWaaIPRggjAUcK
LjIfnDWdN363wrivsLNFXd9YagMWF0MLq1elWQk92dcNijmYJIvI+6wTCPfJBnXfGlvZMR1OIpSX
H65yHfOy8wx4JkVo8N6lhtMFvOoyTF87SG74s4ICzuQXuszvWWi0LjfrWVxut7enfq+0sWuZz7n1
ELKgTSE1sKeXzMYJA7o0BLm7RNWVFdg3+xcvMhx+p7QycEXjchXrjfDqxsLTG8OnsH1Rc9Qhv3gF
CwP5XAQ8fBlMiJPcUfNpAB/O3Nwl+7m7m48wW5e+4XgZNs9P1yu1+LbuUnLJXoBUiBN3EwXzyeSa
qWaURBA8qtW34veOMlOt3zEA7/9EJrsV7jKSOaMxFPU9YyywGCXZMXTmLN8ZXE6a28XzGrkxCdh+
gmW1jmNXOIz20pD0zVBjT9DSGbPzudWvkxRE73NQGfYBORfWM7EYhozR5hFxRlqhYq5fPytElOsW
T8NDQoDYYyQilpXNzXYbyzBVbzQdbUbwVj3lJpWKFJr4J24kGOuF57TTTXmS6LUT0jbjNNJNRbMS
WWFaO5pzNEWWVZPydNlKEZGI4t6OnGT8tA7VRUzDKuyiBeg/j/FY9PKiGUIC2qals8SMfnfepGCe
kZ0z3vRPat4mznm1wIX7rNFJms5V6glW/o74bRPWX3sJHhJgaRYqcCI3514gZ8qA1oV4WlUE/Pgk
Nk/iBstyov8ky1HXrWsmy614+5J4SR/NZGbKAL9JdUQMwrnM2DvGJfP+IWZSviOI5v8n7Fx58e/0
XXHTr4pV5oXm1MKIPkVHbm/eXlrBK+0YxzykR7fDFUylE3+w3OdwTv2sjrm4u7xQr2B9W9dTEmkp
kKtovVJVO9m8yiIB584UuPGlZrHCBeihkqqATc6BKvyT1ivuhDuPLTFnEtZqNUrFhQ83km676qIo
h7lyIUyQub6fUqIBnwODXbuSZh85VWtPcFPsNtlhmPy1U0X3bcAQIEd4Bxj0iBwGhvVqguYEtaUS
V0yvYru1o3HtFWI7hZP2UJrW6kxlb4l77Tiip2wuL2qvIBCeJHoOn5pc8XJyaJXJXZT0W+9jY+NT
NxJJP63vpJ1+FSe7QfkYp5G6IYeG/FSRo197BWyogQIK+uk0OzBBzkgOjG5ig+GTC2jdZ/dmRzTg
xQFhT63anmnbt/qBgRIAimy6z3fpCoxDoOgp8kbrMGP4az6D6F2/TzOa9J3w6qMkbVq38UpRlmWA
USyFNlSXB1LkmEK0Yzf4miv3WdizG1XKtY88aCCUsweiklzLLfSXnSgvVwEkX6OSi6pYG3Leml0X
Zl7HYqa84IFoOirkY3B8EbifvDmNNQFb7YgmM5QGGad80qFH+uXZOsrjqGJkTxfqj3X4FDTmj/yV
dPe52NfeLb2k2NjXEUtgEcS9Mrnwkd+LrND3ILpVzfC6olCRf21ax+1yfK/jO3a/yeK/cfOgACKy
w25Bbk3DMyjrULxha0Ig94RHr/wYwIVslw9kcw5oFkwylfe04sNJw585mqo3lwpBriYLG9LBDvhS
j9/GkZIs2b8anXlDCa0f0bcFn+TqRenQZZeotfpTs0xO2tOChMnZ12pzQB/+jhEYBKOZmY836pQe
1wkEnZQHZksb5lt/SMfYXcj0HXlrmFZ2OP//TVHd7sYeUerUvU8CL1tEF1dZsjJYHGAP5j6g1he6
lD+XQx5V0YvGMMSxtvKwnowWE6k9VlmbUrjvodIQRbIw7q90Yk1iHVtO6OwtAKT+mrxON3cEvPlU
TeTtcFP5cfnFCfZZcKURkvvKx7rfnNvPoAi2Wxb7i0I7Ey8dQpjKrqi1g9peGUEumllxg43G0It+
fwtM78JBg9tcIgPC2yFbN1T1xHB2sIKIEFVxRdqxSd1Bvx0z7+LMu/hYdTuzbJfX2EfX7Gb8TLwD
2dsvj7y+ai48dyLSctP6FgplMeiptPg2Bgh4dcMu4AvVOR4LxwCcHZPPZe+XPmBHXwXHXV0SfQ/g
zP+1kZM8kM+bvzagjeD1qG1GYUFc8ScqhTaXXkl0mm+pG0I6wtfRKBmWT+Ze4+9anfFIt8V+CmWr
KyB07jFoC1fpMRL+XzPUAMmUOq3QPsI6ccPZ0M4juKYw+bPeZlICcZJjuoI1GDLJon57nVOi+rJM
s2YyaND2j1iq0oxLAie/8SWhQjXPV17H1Nx01dHpcz0ATYkJ64AlY+okn52ZZOF5e/lxbV3uC0kh
8BfShXXcyVlyVmQGNehDBZlk/6KOF1+xhCWZ3phvyO0aMa4V00Y7e4rMNmiv3bk1FpgknkeOrCtF
AFYDk9TmOab5U8DxKIWjZajmzGg244ANB1P5isC+sMCm5HCQc9q0q490+Rp8/8nRbfS0g6zV3IIT
4aAMcyZ1O0K0XNxXbpBXwBHn/t50ePnuZbKLeeucoHcLugyDhdu1tkKJvB01BIFnj7XLnc6PiRdG
co2YYaWtRIvJr5PU7eUteseehF4Vj7AaqUVtIC+2djIQFx4iux7rQrjl0KOtU2hcNxsW1+bxUCVl
dDnZc00+kEqJUdNaKZltfdW2p4SCSGe9G+o+Pv5fwYLudJA2ArXIpLdp/u3zE6LJkU4eaXcTZ1oi
ObeaK2AlkAurTGXow/VlUe4CRGgZmXXfUADgCWNcuev+jDiSHHxwr1csqytA9qOdPPLBdYaTaCTr
Wwy3TQrlW+FV2ZDbvZPXzqsMpvwP32QQOkVH+OVfdO6CqKW8H5TssGr5Pv4bvIIp/7XzEObgzyWh
PBariXBzAJ6hmCiGUZVQTTnZwCS4FyYvnGPAm38citAkKCeeE3fZHj/xjB2aD0mfOHaeS/uoHoXN
3xDaSIeYAxgn0Astg00ifBrGYJhCQWGz2vjbQ4kTIDPHdeT7PvyrGGfI6AheuV1uG5Tgq1VEU24v
TbeRq+/ptDQnmxO69+2alpq1dpmHkmZb4zFaZ4+DRpLzix7M7bv8OnyylGLLwARePu1flrKZ3B8X
cKyoUo9HGKtkFlKimShGp0JvRl+E64yU1imXomr0ely3bguv6jaNgG/tC2nq472NMKawAEgb8GRC
N6k/jyENZOKxOcv8HY6QYci6Sr9xL8lVow7SxsdaHQPLtl+cybW1QCnH0ebGlMhNvUeGrd+aPLpI
IYPE0DddwkM5GHAXDyoL+nIdACppkj7A1og4t12FPu//nFEkQcmkfXHB1J3Fb+cT0qlehS/21EQF
HKzLitRtlm1UdAg5IRkFzjjrEWrQiE/+tK6GWQzzxjhhUe0SMIkvMEH8V5VxjMC+eVMOyPdR39j6
R8hMAS4nH+RWImvaCercjJWZr41U1VimytXRiNhZ0PeKDoOwNrE6vci8tcunKbROzBlSECLZPSuE
ZtBAypLyc3Eey/GCMuaxxFrFYYf9ctoA0Vlbj54Bilf3QigefC7gLHm6SypCSTwerScQ8ckXav5I
/j1wTTdaYvyP1yjDgeaiCoIs9W9jPuMVhKHciObI/vySD5kkO8J5Gi4YFnNoAagVcsIoLp3OrZEr
JKO603IJn7hjbx3E1DlTE2iACVOACdN/kAGJ97KJx1b0CTP6ijYJw8h53wTc+3L1liPx+p1OA2JF
rT9v4nQ2+CCqWoYsRin1BiZZkE6O5f16a/ZiO4ktUIAqkc4B2Bwyfp3lyMHTvZV78BE729LBBuvV
09rrVvYK3B7YoDEZ7PJEIP+xzP3k7GsvhVELLA6T0AwiDLdqZnym8eJYlAG2YUJ0FHf18iPGe79J
6aoUiR9f/Pje0HtufnMUeQE6TqRBf4ZkmMO3tdDaSz9+cU9aCUn+rtoPwvF8O6SeAvx0OoG5zjAU
651lDl32sV2ESCW1MySOKPZqBApSwqmZmxHPN45miUVlrdEAbUJ+X1eGYHtrq7lHZyZ3/5fYSc2/
WZl2HqWuQAoUEvO2RfS+d6t0Vr4MZ88NPON8N3hZvXQkUPAqjMhbQF82VpdgmE2wkM/r1jMdLrJx
OgVt6imuhDRWQUXOcu2rfhaaDa3YOcdUXOtsP0ix4QlfP63+jakfp6y9hDi0wWLMY+CxAR1F2KIH
f3mBJOuKi1Hrb3F3eU7E32Z1NI07yOfiezF8+knraHa5iwke6fCxwl8t7ehtxz0pcQpcShtrfAcE
v5xbg+8aowwQCKl0CrZw3oMveRYomLKXZ6iIXWrmgc4STCvmTVrtsGU3Umg2XQczhZRKYIwBCkCu
NLu03YQfsDVvaABWHaKbhhEaYqf0kXGrtqU/Zn3+V6efBo7R7B1RwPO973pWjWM0kPvhvEiKsR+h
HQrmd4yQeQ3ERGCzoe2fgp+6tIfMLRwTJD3nWVBHHv5qdo4fvbPhB/9Vqx3O7O1/hSWiP5w5ww+i
y/mLmx5sqOPt4TrQoRonjR1/ot7pfzwP/0hLLwlGWu6f/AiGKQIvYB0wRM3ElK01T5QCbKBTtGuL
UskzM5FcyDcpAOwuZrDKpTE+DSini5M/MqmTZPqdj0s7LM3krRK13ED7sB1HWb/vV3bMFCNu+ixa
0Gte+egaGwMLZ5NqeRO50eBd+TFel5LqRr/mGpBX+/HdvyIO1DkaVijsLTK0ymD7rimx9XsvTLOJ
YdJa6M1k4SmdUUOzD8s/IJi6G4RIHj3d9MTLRf536bWH9a+fSuWIeZuozGbfbum5lE8LLKch+exm
d5DPzNpa+6LoAVmK9aD3E5Mv1rk9wM2VD9Y3JQOF14meImYdQIBfRC6jljPJveotiInOBmBOLsCx
ce/IeSccZ7Z+dM3d3iEKl4kuWIqGDxEMMmPn7lUxmHuY4Ogm3wl4n1mJlGOmpsHAcu5t23U2AUjk
dDAKUl4d1ooQF1nuO+mXVEk/dGBGI9e9xaXSDnCB+qsE8gC7MuQnjdcBDwkkJXvv4UK90/ofYob5
qT+YmD5WKM7g2J2QbXfvb++ZOoUgnbFRZ3exC2X5X7wSKvIHBaqbP+GXob14qoNTKCY3awQvbneb
C/WsjLPv+VVbMYDX4sQguIDRhDbkjGXl54aviA0NFAKbIUxBXFrpdApZTUGpN3t9mH0pR1sDiZyN
+AGM27meG/feqPeNQOePcXc3oh5Se0dBQjbue0cRKRJ/PhZJieanW5HXb4LDZXzeB1CIztlz4AzU
13ZPDtB45MxWL5GPjM5KT7NQu9b5Q1nl/8L0KF2e9bvTVNz06ooZYkiiFtOFyGsurShIy8ELSHB5
mwI/YzMtlpSYuJgZEpT+DbVgbSfZwifpH9m+glQVWgpadRN1sXmi7e7OiW9OVSC+yPKzXkvFLWCO
4KQFuUHewCGNQHpfoRcMXwu0MdzyzSnTHJkpln7MUAtQ4ISJXVUfzcWZjlT5xjTvYQoh5i3KgjnE
YpTO1ufeYBLwWaGGn2pLFnDmM6FL9jheVpAZ72h5kL7BZRxe3wiZhrxQ9Dvjl0AtQUKcb3f5JJkc
jgaoQxuWetw3RCzdpw7BuTHFeNg1A8f0TtQb9vAZHne5JmBBC7RZYmNx0PkUwSs3RRto4hKY1zlA
rasdGYw7J9QGEG0+yMvErzFF8jJiG0ybdt/SeU4eOhcyifNshuaTR+QvNl+A+AAK7QZkC7I/n1c/
i/7gukaALZf4VVo7JTnhHr7br39OesvbQex7U3xF/+tn0SZd/DXZ1gBz40DCc+3vHpIAierMHSqd
FM1wfL4whAhS904Au2uOoNjVjnO0x9kmzMG2SABLsPi7uvA1bZoI0mfogl1GpHzoskHbl2Fusu57
3d6k44jrWPXl4+5M86pwMEyuYfpHNDMgPaf0c8OxTfbmb0gDm0HlhNEX2PtRdufIN1IQnQJpwmh0
aYMUZS6YxTWAwYOdr/0Xu7w2+MQ1l/aeQn9LwKuMYfBXszIErK5g/fe8cfebIyLTqd5wlasZiM0p
DR5IFVuTYMAOcmw/6YO+wLTJL4DkGhs5v96FYved2BZDUUlArwDgMc/i1L7t4aKnpVP8gxBM75RG
1dfEsw7qI4oa6tLZgcGg6eJwwmEP4emGrvXGTs+p+Ig5UQw9jgr//DSt8fOVYgWu2p13pfB+eYVo
m3X/O5FSo+r9l3xX9X3VwEH1g3vdEitpsyZZUjgon0uiP45AI4XXJZd98xCukxSGtxzhtTVfol1n
VPPtLy6nn7zTEtFzXa4RERLmaS80MJN4MzKUYOk6YayxjQhitsW6kyGbR6ITy8V89Ex6XpgEaMA+
EFnwhw01c4EuLFYdelS3MjrOaRPmerlfBXGkW6ibW4M3ZgSclFM4GRJpUNKi8BNhqgn8YtttXXb9
oSMfB9Y/xzKy6XshHPvvWVcA2MvFWjJdD+1v6ScKJTcokpfcyctDs8hA9Emg1b6TOixWPOfvCk1Q
UH1QvOdseIXQxidbEPJqfCq1VHPc+sJ9+V/P3LRw8ydY79825C6Om2FovryEx0BogLHwWl1w0X9L
I7UDPzP1/ppqE4QlnKM72cZON8msoPxekDkVzu9jB3+LoOpHmro5UUN6MgTdHopT3yFiz5FdUERF
ThluB4oQGpFEDafQXm2gRpfoTVzaIfY0Fpv7IXOFHWVcfBWVltEsuQJJ5I26AbIqzpMSqbWL8Nqp
jQKUZBzLzxyrZlmnKHy7MFwFgz6UEw2Wq0rewydlSJ4g428SRPHfn3rLM646ergyfpoZUCk5PQ0k
3+7uNhI7RycGGZAdYvYxFkqa+D/hTmAbSKJkgvVbidGa285/kAmsaxOLZsjNvfenIv+5JKPOH8wz
To+Zd6V+Zj1rhfLbkGgyldqN9nM61m1OGpZRa1vDPms85ingu1cy8httV5Lf5gm1WF1t8opCn6HP
bx238pYw8nk/KK/H/a+5EF3WOYe0u/cz1FPXADI3zSljiD3or4xF5eVb8oHVd86i/cMvJD56UZFn
nRq6dcj53XVhYVaTtdjDGz0O7ibJXgtg/g/DOAuCCdZHYxzf/IV+vStB0879eN57PbwqCXsrJHml
z902DsH+rLEoOatTMi3sfbXHFlIxD+Ef/i8qIjh+FhCOFRpeU1AO+ZVtgsXXsqRGrpaPgykGD7nP
gEssFNO4br+Z7eK/LY912nO1gysoEHbv2aPUyvqsXFuytrxi6DH1IsfQW86h2j9x312iVWs4jKYP
Y8+KkftlWybnCArrBpV7a+4upaOQDN/Cln0QVe+VQFwazV8nXmTnrSUBlW2gDvY+tJPgv3xBO9Bl
dfpmaBw8vgiURp6F2ruG4muyEDfXV/w7sMyjiqs44u5voBQjZymHDxn7JpPsACD2RZd/umshDoPE
bsfNbVkgfDI9H2mEV3z7ts3zziPvlb1fA2wbSBRA3R2nCMLsBtR/HDY2u970nfQlMwRRhafgg2Eq
u7PLUhtW+bLxcm0mWboR7JXHeTWmj6nW2c2kxuFMWg3uq+691Q4nJSsEGL/mqh+3T7kRVJfmWmyS
RuBwKjuLbB9/XKc+DQzf9v9HB11Vc+j+4JE+JVOd/ld4fqWdAa6WaJ3eu9SgeYcaod8DKYuz5TIU
EymLNWKQScsVqYUh5nf/++tDJOptejjYLnTSHH76igV1+yqnsEEvNkd1drR50yZo8wrAPJj+XP4n
iaqkGDAJtfB7eBe+5fijLJ+T0R+fI8qkvQGZi29/NppyOUMcn2ZySsmLqjHPOll701B79nj7QUf8
KJJ+la+Rjw0TC0k4QN72w6b+mWMFwd1+rV9fY2PAzjcnMWLOb9hknvBmXvPVV3YdGVHf9tNEpPCM
O1le4lXUmmXzRBJM0o+fcoeRZiIgjgZrWrfnLHIJ3LJfmay4Od3EYcQnf653/wfVMIG+59WkiyBu
ph1CPUfguPoD7HGH8cnhdNYcHlevjF1e3pP7E3tMdCPHqkmyovNRfy4khDhuSnGGgZylwju6yIXJ
3R3oNmhuJSGUxrdrTtcnO+YD7/+ly3FyofaoWMEvdjOefhKw46vw3fH3bRNEcJZA8eBSH7J2xw3G
8kki8ETfiB+camC+ltmMI9jtVKJW6Xk+kKcMBvB7oOqYjmQy/H72ZaPQn2vcJM/JiMpe+PYHnIhG
wlyiF9R6cccMdUghlRz6mwiU1c5IkYr5gqbzgP0CEy3ceHngKKq9+5NoLCeaRNlHZIiaDWCO5lJ0
MHgJOvX6X5EWglM5bCtiNZHA4tbZufURBE4JylgUOg2uMSDVES2Iio29nWnR0weA5XfZRUUmXnK0
DCHEP7vQCMNTgSq8Kp+lbELEXTjS9++k1pvloEXbaUywktQmjQiinPqOzXK17wR1ohPO9ghcc/1u
xYe1pindkyto5k22HGRQeElZeNo0Mpd95BgTXblL1yDBPfQXtZG7aCmBuY6QMA0T4c0pcwWLYYO5
OBtSbLcB2USwNxjm7Dd6EFRfp7Ge8NqUffuoIz/d34uyNzzZaq+57lJ/6jAXmFbySpUz687J2KxB
NkKPvv2Y5+74SJYbrmCYOTx56GTT7xM6o16syeLqnhdCJogA5HVxNIi6qKyyFFy5cnDGmS1Pvfff
boPyBjHoIcENhrmIBjcwdBoxu29YsRHuWeruaqPD3iVzfPs5S0DetnuSLyOAI6alCsdaImqsFsqR
xRMykUnsw22nQAh11T3iEeJIlmw9QS2xZufrtGK3RVEJE39x1eSiiN4lzasucyNqarS7rKSPaz2x
N6sDv/DzWFERM+sMGrF/ZvYWIIl55VH/zAOb6P+ZTGF2bFemDXNgVGa8GDzrc1+DpsmnhG6a/gv/
rbhapYBeGAABENkBqZ2zJ9stcM0wrou7R6hG680xtI8XEqXXqn1AS5T6qCQ0oXpfgPr2BKxhAzJM
DCzST+3Hsqjlpot4ywKAWtEPybenG1oKUwq252+o/op48RUxtiHRGIboKq4FpYl++7wfehbc3MD4
jsU6WnAv9Ws/ZsKf5yr073rLRXm8NYN3DlWvo4W0cffTgFx9VnB8y3HeOiBmEXxbKaM2HzBje0Lz
6solZp3NF5dDN19MPW0kyUzE+rSOmC9WN9n0vFHHYbuySf3jaqM/Fy2kXhzIZVux/zuXNLsgPdHO
4zP6eeR3TP3FmFMc+3Akd+SUdabCbNlMe/+cNtJJp+I8FDmurkpVpitYjIyhOySE3a4tN69ViXVy
jKyl4S+hGwJs8d1KisuppKlA/SHIk2nENWxIsD6Fh/QOOd5FCDH+S6kTXNXKeKrY7CDf9Du6Cv6y
gFEYZgDICi226zhIRs3GkWgXhRvLT92GJ8pBkHd/KBHP/xpjbLsF/I4UpEI0YWKRvDYgHSAFOk4E
bxVzmqYUljG1edYpvnGVecX9c+hO9hYRGbA/UDgTBvxV6pSjy01yh+z1U4qFkZKTpZ9mNDjgTM1I
wpZBTcvQLImoxd2WsmgKiEN+we8l40iOI8xmrGgstzHtlZtBtVp0tfpKxXmC4y4FTTem8W1m8+ct
+GToT0GKEWfRZC4atiQxP8KsgipwyC/aJf78pnZNMck1mUJrFUIvaFQ0CEwbyG1k2ws8/Dhvtnj5
T67FavqLSEelW7YoX4UvZUuOkn0+A6M4pgEKUjAMlsMh/k85q3t3BmVUi+QZR3BekV1m6fDNFYzt
QnpcyhKj1845AJnGKsXWjN38gxeA9/LWM0IVcjmwn9tTSbk1B3kqnAiTFL53YLSczjIbVi9wi+2B
69EsTpoU24p+t/XDbjwgqKl37mi1F01qnIqvxXCmRblut4SlPOT5Zy08pl4ReRvO71z/I10/Z347
HfhiglD0KNrYzx4UEkxjkmI7oJVRKKHvYNjtGpxaZ4UupIWLaQYHeK8V1yhITBZx/nUiWZ54kVGL
S/fSIPQ3zIIGaSDrqaDJ9Nm6KmH192YwXcpR2pXzhHj79eMYoPTwDPbtonBNRz5j0yHtuoeo5Pcl
iv58t0o7+J9dQTQ65U992MOLTRbBQkk/ZSBt9xaW4JgUNKwAXp1o1YyDVVU4Woepk8UvfTF9sGam
LIQ7jICl2rsm0Bl5foliSm00X7TBdrYwPSZDgg9s+DejnyWXxOoHD7KvGev7TuSkI5fnkJBL2kPz
tSWSGwCHe1S25Iu1i0uUJoF9XxKBRsJOfLzePwtcbXvlNfUHeGGuvkKlbS/W1HaYHoxx4guHKxNV
x0MSZI7kjiwSILmn4APyrtit+RgO9JDY/hep9GnBMrQdwKyhNkrG8AOVW2e52OXWntBrR6VLZIdp
MORjR9+STnjlvzBR+5dg2JxxYqGv17cYSQ9Q8JKIkCTRArav/P791yX37f+3+72n385j2dPNGeUn
jjFtv9mTPDADQdd7vlByjbDowCjeEE8RChmKHauZ2Q2Pt9ZcXE3vtT2f6qiSMjN0DI5H9pQh9ut+
Sk9xUPnoWxcF47HgvJPVyZ1YGw8plwHBGu9I/D6lZpyIVuYH5c8QFmDPYutUlJYtvvranWKXwSUM
OvF0KIhzIA7LDo0ovYvnOvnz8c2eBpW9Z/12RLr4XaYWFSB/aR3G6HM3aAq7pW6BSf5HbQ1pR63K
mrqvstB85QAtPE+YQUMWrPyGjjQ2pyDqdnMuPFdFvsXXxBH/wYJkZiSC9z6Kt1fqMt2vVTWrD37f
jzwM8NZIbj3ObRrkrHYX4qoTbmnZmOkiCYj6AlORQJSDXkwrzptzkF4GHJlg/5d8nGUuWAjNao4f
UhGq9E9By/G/0wMRTcI64TRskB35T8qPTbZ8FyJCAG/cnerjPsSOe1QsWVVE2TVgELpW5L3Z+Cjj
TJ2GXuLe74tLkQ/sTRKoJVciVPCuTRrFddq0PXRfmYJ7QeM7TQGWvK+YygxImeIzZeIZQRh1a9NW
1BdPKSaFYMBIwSXQelmHLukiOqHyVMcii6J9Pf6UJFXBkIu0T3ASF/gL1NmXDiWdq61l2ncW15l1
WgMy1WbigJdv7xwiqbW1aeE1vJRxr/l85wbbTqS8iVivONwNWxlkrOTAGUKU1zcib618jt6EhHXK
pZ5UgvUNEiRwd2oNRAgObGO7jRF5UzbaaE1TGyoE7s6wzOeSKQ2OOfTLBYS+7kGKnKcxTApGcDnZ
U9EgZn5Uk5ONOv91H0gzBhDgCR3BlbVF1Mm5GW12PHno/OePNgGORMxiqfReas3om1VHeiSee/NV
skg9nQGMcxQLDYJwevNxUZrR2O26WmZpbFoXKCSR5nShz5xNarvZ9CkGHsTYG06kHWqtNOexjsip
QQqez7Nu9Y4ucmtk/cESE8y3ZoS2CXb6EfobqzaOWoO/qI8qsN2iSNP6SHV3PfVpBcQAxWVmpvNX
8AXAsaScPE+frF1PG/8iuURJpdb3TzO+bu4nOr0u+lSs7usvWvHSAUeJN56S/55PAHFVhTrYBOOz
9pe1m2Wk92Mr5QO1NBFdSeWO1nQDEEU0cl0lBIHx1PNz9uChCh+lpLq4ryr/0NLsbLGaGmNHHM9T
dmZsI72NuWZEFVHooF7iTkPdI8LfuUT48XrimlvIUy1erWybCuD3k6levqwhNCHYG14L9c46ff1Z
AHWPKJJxoYBCQjxF9Q6kC8SDBNk5sGjkMJOS0Esc7wNX8eiEoXBEFdZDpzZvdhaVnniZPeLRGAO6
DmG6ynqP8R5jbVYVYXpTV1jr+UbYZlGk3KDdwz57qcxJQL8VinL4zxOlg/NZjtku+AvqhsECFW02
QdVxyegISgBP5GcHOrPfy3+d0SKUsjHJ6WgJusXuXblO1x1e7F1UZU8tk3M8jrBEp0wyIi+TRneo
3wlJ82SyhaWDvjz9Il+54CF+f9ZQXEvVBlPsVduY67z2FSaQZqiaEC2DQVds1QGe2uNqu7wSAV2i
S9w9VZkwcD2RfjDktCE22CFKFoMc9o3FMo1xM9J+FcoDJtxMobuUo3oVTLt4FHzVvGFlQBzzjBT9
3LOcWu/gfn8mtYDvun2BoxKEOQ1n8PX8UuayDOqsp53wmNG2bC2YEUVsUmQi/neNu3Vtu1esPsEK
GCMnbagC7bE6U426F0qo/8RaKbtMDLOb9jlblBq5BkWNEN/+lg5Zer708jSk6t4dACvfyM3bFbQL
nESyfm56G7hcIFfc8WstsaGdjqg3Qw8bynl7cdh3DRRInBYt0119j3uS2bed8Tgb7sl4OHl9uV/w
vFi4Ho9z3rcOdsCGy3KdL0ZcBj1AjWI8T2mCohFvVoocjZW4uY6GFi0BdbyE/j75rFsfyBWwvgTV
jutu5XjAKAu/7nIQzHY55dZfsCbNrZYFH2NlDeHOloA9fNcc16HsIA7GcSTJkj6gqFG/XE5vslJ+
7/DrxVWs/HFdgwwfKGqemCSAvYgUUW9kiD2OGryjFcFoBFxIXuzQYYTx9brmY5zwCWDVOmuY1zLx
csL3SyEn5yxRMXWpkdYozTphJDT46FXsdcF2xBaPN2nqVzu0UDv9Ht5yzUvonEQLv9JJJ1V4NEMW
Z12XXL1XpoZ7fO0GT5qX4h/SjPHf1lGQfR5PRihhlrkGBNjgQh1Y5ssIecETE81VzUt64eRRn2Mk
rXWra5cOE4H1QEpz39+N+B/uXED0Q2V3XbqdkQDcKJVOVaYg2qOOlnsZzmOuY2Q7W1IxkFmPnu3+
5c0y3uhZQeTgHvKRj1u5Y2W0Mw+tf6q+1RTo56B1zTWaXv4tvTPAmLlT68YK3Y96QJEcm+tRx59v
Q8uk8EobiRF+fnCixhDkIF8XOexlHazHftlfBaUAQmhGG+ikQJbxS3RXPJeU/7X169Z52qvLXI7f
8l9biJMl5SJ4+zkmG+hqjXgXsf2o5mkJaqNiQjfoNlsuHj++tJawXBaP+P//ka96c73kIkNUUQsP
Kh9bKm0YjFRO6VdkpANIz9HKFGaRwrEU7Jn9Sfgdi1E4toPVYWe6bMZzSOpvDh0r5I8dpESOvk2r
3FRlX7kf1BX9fHVWqlnWw4197blqHCxDqb6mPeAqOntpQrHcsHe2804xaPx/uoZ6Mw6NyGartDCr
1dW4OSjFxOBH1r3u9FKkt/AUf98RXPAWOInnklo/qKNACndI2Iam92zYfIIumL98dNsCGgXN9kBT
axBNnvzhcrU2BmsZ7ds2/Z1CgKpxnoHppxoKBEjoyNNND3/qvSON6caxIWRrTC8z/8DUY/GFC6ts
zapbU1scJ8rHHWDeDJohlMR+ePP3QtaNc+BFE6OXwFYNUEpelImD2+mcs+Ztl8oXZWd2i/1nf76r
XqVuOZE+88kmSItzNa16+OKfV858OB8zfwx1VbEhLc0/FcCN+LSu398OmgZGRGEb0BpSRqm0eheM
DFppohWxhvF6VvmNJvqIaerdc60DARtYCpNPIWssKFQkU9B/v7ouy/p7BQiEw9Mlq7dCuhPHHEfZ
XzQ9eVafwN84NkoUgzuae0qHlQMWrdak6KAjExryML99KZyKW7gk3BG9FB38DaRVpjhzRIpFdJol
h92166uQjUcRI18SOQ47s7jL0z5S70AezeEHQjsdrCLU4bn64HynYUKfA9nl8Sxt81Hv1etjHJ0h
3HPa8CkLgK4O6oggvkPRTuC6pTTGePTbIthSHSuOKmYzxdkxpCU7hxAJm5MR3wuMysDvtRk3fzvh
BLPj4q3K0Tt0gpbjIINNSPv2sIiJqBlms6D1uGE6q1hx8rJa6t39KLsBPCpHwmXMujLTGyhDHe28
z9C4IICbSs6aCRnm7lGrbId+hteJckgyRg6pVd0pOp405sVPOcSUPlUkxmDLiWZeP9cDbYkUktLA
5FaQu4XsWOpcZpmpgizX9ho877Z1xp+zvAjAaWBftnTmc+SpVHi4C/t6ZstJbsbMiCLGDiIpKFMm
FaFUuIrW3ASgM4k+MHXaBzBNT18k2DbZdDzl5d0D6LR7IFMZhFYq6Ch5+bXtAdGKGy29o5mVVbXf
t6iQxk0iyfmeWw8Fv0LqaKZxtEPJMguxJYGDoAwQjCPvmxzjMpTr5WnG3IPAjBImTqQIfJ52hNDh
qO8jYTLRiEUXlhwmFETJQMb8+OvsHY42kYvx+JAPqTlY5ygoTA69b8HNQAYhlryneekMqi8UbwRG
y+fTD9fysgLMe4oXS2nAbtik8QAEPqhZNxiudOuWgUuuY1fLcP8nyCj7SInCG2mWs0z0Ll8afFRw
OjWYt903VE9/5cfoWbTd33ayR1u7qCvLW1ahhfvKYM6azh2dD7TTAZ+UbQWYMHhl3KNNQ82U853m
6Z+UBb2sRSS1f+pnkJxunirF7LKFl2NC+w7dLhM4DJx7ul4m6VNXzPuRfIjtXfy36OJ7/BVe4xmF
7M+gdhYB7S9WgrS+rEOxYcYLoRVr2pveJpj+JWZvL+mIaQajJdOU1cDphXYfj8CMN3TgogIDpAFU
IYQlTau0c1q+DUQnuKsXU+SofMSO0EL/+NwEHB82W2vbragjdZpGR6SocHLAJfVyjW7d42rnYOi9
XT7JcIMnFjtSMP4EK4JeTUOCUUJlS2Ab20nPULVpB/PbPggrQT7NBWzVVj/BvW//4hhmT9bdkuqA
N7b4E1f7Lt43FEDZMM7R+QbK65QguWKzEHHEjvWv/EuvMqDVnTI6vYzFd29hWgn82e/DNgvtU4Kd
n5Uta9AttJZNkKkd+T+2ge9WuBylP4Edjz8THCQD2MwkRgYm6Xxs1FSZvbjVco4YLTCr8u8cxnm3
JmLa9JAy6FJMrwGdHcv4xuhj9Qo9Uwu6iWT1lMNcoINBWPM4cVbiQ1JgNLpuGckxIhnxZQJo5YoE
iSTDM+6WOHjmfG95ZkeJg4V6dFr9evPAuWUQdXvKop+V3OMnRWr5joTYmHha0jGUV7L5IWariFTG
xXbH6ruBYYTO+NBGm9Kk0Z8FVVOuMZRewl8m/RuYzyKOGfkpOupJif6zvinHywwCZY2QizNdzvwS
EfYB5ggPkFElob+6DgX0aWZ99YGDPWoCRh+Pir24YZ/+hJbvicSxlRT6xkzXOatrGDFCDiY6VKjM
c/ZhjjzSNelPYrpstCPQkzqp4vDI/4p6UvcSdT64XskeBq0eMxHmwULJ6bMc5+O9S1iGEjRkSQtm
gpzho+7GGbckO+lkYZl3bnQZh2iVIEWgBwvHLnPuOM5pyRHYOhjHZtc551wauG0+JuRYBTDUXo7L
Qi+o1QXB5go1M3i5gSigtQXX15n0yglRKr/G8JBDrbMh53Hofj+tx5fsd8mhaRuQF8fcH61apoRB
BaZ0y+BMGPPOX6rGt8Wa7DMo6RJTIM9C5LCsA5dx/xxWXZTBiUpPPrusfGvUGApDt048ErzKLYlT
OthbBAMV65KOJKstj558WN8PN5EHqRG5A7rkPKBjzxSA1sQ/mffvGzkIFUErYmwDH5Nr/q3Fg4Gt
0e5kxaqZmjgolDCwXVFT1OuBid4/ICuTmXK5NhQMYVXVwGGcVRyQD1n618s6FWh5pMy10WFUfqlM
FHBeLyau0Li+SW+ymI1vKvb/AtqktXuvSiFiUOO5rrjeTkQzcPtuRD9L4AepdH86EVAg8mLhnZpl
zOKKXfrz04rp59nBSFtSw9m6pcbP60vIGxcjeE4RetwgdJnDxjQD2VGO4vMpJQdsSqNeOBrJatJO
yM5rDahY6Yi65m+9u75JCjTRxNN0HI4j92KWqu2Q79WAO+7doB0zcprnCNHxHBC7tQa0RapFboYR
FBf8HgN6j/61ptfuz01ViboU1FfQpJftwFGwgRjmJepRzmSIodkFieCDxXA5qXHxe4JTwEKSVZaG
g7Cv16pSobeTq8v6zd77x8R0TqioNhlW9p9O/sC++i0zhUZ+Wunj893DRXK0i+vDpFVruLz46MPU
NOqCOrs2mzSuYjUU0B3+zx4fYrLw9Pz1AEC2Sy8XCkezdXGYcTBo9ETrPvvWf/dv7R1zchL+Ivzc
wf4BzoHOWraWIDNf1quBt8lxEMhALLrrOwM4bMa0A/rXcYznffdcFvVCWlR5lXs4cw2dFd/OhPFH
GpqDSBHvCqYad/WOlPR9kDG8JIhGmy916TMIm54xh8+zsSRZocoZ6SdjiVJJmG6KtqNRgN2+nEAh
nvGlWTcc9WKpshThMIbRjtqnhDVUnoC1Yi6rSbbznJckFV6etEkEP74g8pjVXJ0eR9xt9m7MnPux
z644l7LhsWOESlNtnMPgJFKcXvNPNum17fU4v5mYrC1V6uSJhSUV30JEvdzqjSx176lohyHIURVD
bi/cESif/xaX7ae2yQPMAppttNMlhERiiT5ifT/qohjuuWKTyLAAy2TV8x618PR3ABoqXRrANZjC
1T3RBVlw8pV5lhm01qpqDYyDxBc5nKZsyHsQcXSPhClMOsdN83YmWmDnEPS08GXUFVInnCRLvm/2
ev6CmV+usfDhi5tL+ARHpiFDktULnz6xSGdezSp7tEarmJUmXj2URHXTHU3pDtTn38EaZy6bxUFP
VwlC7A3dI26UwM7XmWN650TCRKoC8AzXr3qGJvIGWTORQWUG4RicKq3mulKmlDNLvZyLJ1XUfB5H
yolfy1l2qb5loxn0knS1qvq+BiuNZOEx+MeokFLAmF5N4QfEpayM90rseS20NkWY3hDJ98gArOR6
eapHl767ytDrpMjykdHVmGS2if/eOg4jUsamsQz8ZqaYNuFuDtlYn4f3S4boEDPwf6SYGcxxGiGq
kMyL88S5QcxVJlm1yZo34lgPPbd+c9+z9FTq5E2bEYNz/hZSRcI8gsvaMNbvdZYZqa3qf8ilMnpg
lCHviIHxap9WnVFmL30g42L4/hWtecAq+P2YLkSeUV4VdzP843y3fCvw8y7qU5gDRdV5lgE+aCB2
dzc15oOZZwUfbuivWRSdE+iRmvxRZEbyMKuyoPoe77H8zjnHIoDlvq2GrVx1jAfTmQ6f89BgOcAM
UiZZJC1QsLwspe8KvhWbK6l7vkwkXfKdSIZeqkw+83e1JYCU7dt8Ghoff9hxaS4DijjZSn+aj07C
Qdep/Pr72b1xu50JgQ26XwJvXf4bf+rkJ7W1srxsYd5vcbATHRV6sM2v8LPMbQMLvbYTMLXdfc/+
OIW83wwTKo1Tn3z5gssmBUtjWuhta9Z/Wei9NBrEl3HEoglX4DRwcrOXxaAhAYZvgglhYtrM7X95
N+jEpblBoPAfF5rxiZNyoJ/MKisoNueMyochz6A1t0ggrKXMXfOZtFqN3zCjmx+Ry0x/GpAfPDdL
MiTG7KjtKv86u6zP5NdZEE+fdN2tIU3dKq8iB/Q8cDQiSJHRyno8DeSb8Bc3eTyY670JUOYRJ9pT
DjiB278H125Dg77In4XLZKFNFPnqU1h4h/NOUaUBohk1IUoTNQz93oEhUlbEOVsOodoPC1fupVMS
Gw6saFPKZanAN26/Zau+7fsaJET/zHwZVV1bdmwsTDvJ8q9AF9YhHEXl0K5veyoGsj7qd/XiyKPJ
LUlqhq5z3rO1iJTj8e8jOgCrNc4aQigeVre3Kb8irc2RqXXeR7AXOxypUM+hgTQFgQHN0fitv4Lg
ZRcT++r8jFDwK2A4BbwBQe3EL+rQ4H1SfhVaWCw7PqFbuXosS0ZFBxNjSp6Zfp49SSmjtCPUeSkH
hlCIJAGByLdWfatZPCOiJkRoD5SRCeUBNSkESD9yD31OyZd97CzMCN8moqXIKKv6RUhiflBTB2yZ
TUyR8Cgh4N8KjDNr88CqUHSfSoffQC/kYQ+dEnwOyc6beKjjvZ9jBFdWohynEb5dZUt/QC2t1Ytq
f0yVOjRpBSjRs5BxXQcpBG3yJJVQpRfz8lAarIjjvKICBpWSWLHrm2tiZGn4k1ZGKYglsTH6sQlQ
ucu+CJ9NPa7KMw8wt6ikR6fZtMc185qU/upP2koFrrmvksTWLZYkxPuzuFTPBywQbw4ON7Y15KnE
aFYxZ+hklZRLpSzBcJDfgvsSaDfo78Dzs5+odpJXA0GqvIVNFjOeXAhh9Cd6D4ADkQNpStoB6PKI
2SGnWyVi7q3OFOvgKoA3PxDGoOFN+ZgYUpDO/bzYYnlh5YCSt5BPXmSG2gj7bnhzzRFn4ijkbHNo
VoELLjl8SqmIaRRdpT73i4gB+l3M1VcpP9yKE2BUSJslfSrUfxkd+fhQOBVDpfxur2zyEHG2FueI
ebZUSSAcCf8ski7NnO8c9MHAq784FWm1NMTRkcbdB/nvwUc4IH68FkCoKcB/HwHCiiSFsx9egRA2
CWQKlR1RrVTdKszwiCFmHhAsfv7Bo+oFPXYOTuLFazynbH6AN4sIsmzZmhT0Z7K8tu1ytFlUpsGK
z+QByOxknyN5q9sftxY509nCclEf3mv0KAZ5ORlv5U+agy0AWO9d7nLtl9jV8jBfxyIhBJoxT+Zo
hXBZk9wnasJjxNZZRmkHEpl/WE5koSERtH+P2l0KlC32iyAlwMuqSuKXlV2vzq9zEqj7RSDOyDKn
RLMzsH8b6Nq3R5xR/AIh0klZParW2uSfeSUQ++wE9e1gnrqLFiN4E4E7PIMwHkClzJwYtRSt2Tlc
4Bnbrd5fE1JdP2kEuR5qyOwq/cmJn8zIlvY/gbs1Oamo1PCjORv1u9eVcpUPLXn+4Nioij02FCfF
z7e8QQIaQlymKNrgNZvRlmjMwJwT2arzepPn+5ciLBGYF75LZ4KJRfXiQzfMKloSxAlyotwKV11g
fr5WDlVsO5LjUuYjk5hgeo4lhRdWWKIhPg8b5ZhzmOTm8yI7ahePvC/JxpjvT523y1dvI8vLrvlA
UvVlnT+qljk66qR7zMC85u54Fwxqxi3TUu8z3qYX5CEKtwD7QkIDB2SmBNHMmPK3+oH77O7rqlER
DqKxPyR8x6l6vHPl3RFCNPmIO+JbB1Q5CP+v9ot3joi06O7ZIZaoidJXHmosV/0qxTteBmchgXF6
PkH1w4JlJnJxpql9hPuLi1pIiLxGKLRZJdxF5/IXcrx7hAgBhA6Lz3hjL4ofYi9WMn/MAQHvuBK4
83oZRwPh+eqC1qncEu4UvRQyHvW+uhCBtD5WIANZ45FK/SWrErU3pmKo17BCm3pGyt6Cl2t8j2np
cYLHQhWoFA+ig1eaOLvNwuneDYnjTz+gy8OYe0oTc3rfgitxri9ee0k7z8a32wwA7jdrvxVFYPA2
Bjq8iySh0lRNLGwKJsU12u4136ydNmdpH9QuB6P+nFgVCO5ZUCwf+5D1YxcCAigqxpD1oEo//N0W
DJqF0Wf8S07tkE3J/vGB2N54xVWsz+CRlzfVmuomYTQDEPELBuRdyqiupS9Lucj/GtwZbVTb6nmw
Dm4Cc2zP8NQ+5vn58gz92aODKtNJC2nFCuJMIX39gmRryP7s9Iuwqk7idfQK29qsC/iJVQ6GBhQ8
XnJhPGKrpGt6IQgpNnhf0cmLGEyAlGxxyS31J4VrdPwrkhW8+IUl4uGQvACPdq2nXU2eji0tbcF9
7QR0AScpTp5/JTeoOW89j++H5xPm96REcueoV9O4i30EEbIE8f+VtL0phG+YZrCV4lB3zjXZ4L0C
35TS75XFz2QgwnLvDbWTiJhYFAK1+EmnWcIwk+RKc4Q0lXfkP1ixmasZoQmFCn22fYIb1ydpPc7k
f03GQ5zSg61nQASA4Vg5I9VLcVZaaYUffI06GdTPSZ+Fq7RJ0ZUacEICRA8ojq0a23UkhBWpRWwW
ZUAerEUZLsAOacj7xTybh00E+rNy8nzerL/VVrX0Ubnyjl9VvOYeTIri5nSAsfC/nlxMhzh6P7nE
xQaaCQ9rKVXPIhAjKq3QDgv3hBtV64XscWFsFtXlre61xt01pcUo6j1/HT/5h8tlwllD1RP77fk+
XmXcDTzz83nlZM6JzNrDmDbSkNSxPo6v/VTFBbilpSVjHe4MDcWTMD7Wz1D2zw14+W1PwFr+xNk2
QMHSTplBGpwtTfHikppmeDIC95M57Di+d0KXBOBpA61fwlIXPB1q+e5wQVWxNxaCXh9Lbj8mIS+U
rku/DyWioS0GJNk2fVjwVtCB6tNj1m538JczhfPfVnCRpjV2pCv+avQVADTLXViLcxpd9DOJdUWx
ALTCMATOslJCSpqelaSb0C40wLnPNaQGv9dIZQP51Y65hjFm20IfTCGTFfbuYGFzrv5Uvlb8DPbR
AEUJLso591fthFMPcX+lKaYSzGFKBm7QwcyRt00aCTaxpwN7vjuchwFcTnzzMu/hJtfeWwEZdgyR
V0b49YFxKtCf3bUhTr6lRow/17nsFUILyPYKb2wx8aG5QVAd5EsTPlDQcrJfUa0PVnIIqvyb5Qsn
P6R+aES0mv8jqKsD2er4fhftxBsWRTh454sT1mXnQ4tZtoh9db8w7FTrhEnFOr7bYjxaBDUgLjj7
t8Srovmco4yagtq8kB9Ghc5fdRmzQo3eK/K7PDngFrLG02noGn/F9I5HWohYb2deHW3w69unoRyA
NsxUdVFyzhX8yZZE/fa6Ks4PcPQ7r8shJ7YiGBnE4zuEgJQqJWREWud1rhDUz3mzoLVGiv5ax1Tn
VIlhUDvofKK7SXw929d8C73iDm6Tq1zX/ixJhxz8+tNfgNmPXgU2yr8r8r6I+Vfn+99soykH+ljK
uh9ATxpJGks0UnVJfQ8nftOWLMIeLwjPlpXzdMiHE+LWqfIaXLcy1IHtcgvTbJb58Q1dnCsaYkZr
fcn9gLYoa620K2yhjSg9fjvaPWXZEjAxxPqL1XGw+ufPQmYhEjaQV71s2f5/R6YN9xp0PBs4geUc
iCXAo7hewDR6+aMYvlV+96+oFqSJ0B6Zo6ogZ+QDo0gbU9pQgWPotcFFTkuZiiPmAovDH7Dg02VV
uYZdB+vAdYc4ihg93ghxz+3oeS02jCRQLmQOfEfAqDc7Oyd/5y7v45DQUTlvBv4lsl3nYkXLaaIZ
f1JJZz0WuP/MPxJutztsTd7hN6rc93Hr9BUrmqYRYf/UD7NgBckxT8nBrW7ZMgW/rlj2UqLoIH19
Sv6RnUX0RD30oS5D+0WVjrmRKrZzcHU5ccH1FcxVk3RC0iAtZImKV8h8kBxzH1FYztmzkUt382J1
Vq7jCr8lhcc70WjTZMesQUEmIdIkFwlZ8i1rK2YD07HMISMSEw9mDolx8qT6FlIeL3EGCUXgCOix
DRLrRujQpHSYQ6v3iDDi0pACcRhMbKv+KuIjsWkB+LO/YtHPniQjyAfcCaSpv6CmeZlgr4Au/lmA
LX7QBDMc7g+jGTzMirF8MznOKhHtkObCi9UmzlVbbASXHqPD+NOCDDnmnPniiLYkT+IOuIdKlAwQ
+S+34WlZBtTrYNuzhVQIiBteVyRmDFcfL4y4sMLZDOjAMjrjstF+tQt5cia7n4I4SAydKgI3EsXQ
SpCXLAAPCfr4uX7djkDb7/CMcVXHsy7CxfZGI3vlYf3XtBTHaiIUKa9ccWu3dB93283dIG+AOJ8N
x5vSjwxduvXUBLbmXCp1A77FTkOqcP8I4hzU4a7/Iv8cMcuo+S/6hWeorahTB2cb6G8TVHqpM/L6
hXBAPdMEczpHf6kzGgtPSCEncKdal51ni5f/LtxKE9PSJY/nui83JKCKWID9Ayw/XltNNxqDFSsU
YBDIA9Zfvj3fAWWU0pBDpzT5//6HoRJ4IS2HkxBLObp+En++2iPNCiC3IsuAW8FCx6u4o+zbY67i
hCw9CQBEz0CPOFz+Gjl4mcXMp1MvRc+j0sUwyWX6K+t5xyvtR5kK+96kXzQ97mBAt6oZtrZiV22v
0yoruOSnj6iAB8awC0YLuae2VO15CmvPsniUde+k7lSiKvOhVE8qCmFQnREBIFA+D37BGHIDCZuP
8iyhvUTM+H/03fcKjvJ20DxsvSGczSO6lY9kxM+XwuVIIfYdz6zv7H4EjFPZDTidYpLoFuCRF2F8
fBdS6qfCcDRTTZnYhOc+SCOjqudeLiv8vPUeE17/xkLNjHNvmhq+zJqcdiZaWM36FUwqOKH/Clkn
gKs4d9DQheuJX1lzeZqUTubnnwwEU811KA4h0B5J8oLs74fbSvshRJXBc5qTCZ21lU3tcMGarWrm
PnIwMPFXrWO27TnfogMbZDwBmdab5pe+6it+OF3DLPMqO1Yh/FTG3Huj0vRrIp0bd12LUGH1ddVw
hIZ4s0AKJLqwLraqPBAaHB/cj/20jDcScGwfuX2yyVJL+/jWUen2eM5PUz/qc4LtU7knjdoXOSZG
TfVnd7uZrcsWDXu7Fv9b91D19RhwOVdoytVxlcM0kR8doX68tiJcGBvrcO6AHPS41hgOkr2CNiGY
gjYRfAXfqTcwO6DFAfuCVIyZScT3vf+vyUXUhRXnlZWT4DH6Ydgp+Eok66oziDiwg+L1ZhrjBmTn
8UxmLp7O1koJJF/wgX8y7KJBbbElFKnKepMKary9C8+tAs5RSUueHKz0eyWsQ4z7NBNj8kbvvpM6
WYlGdt6XelLo+g3cke23yyJTF/z5En/JEtIUeRrd4VAUOAls3zHb7CvUiu25+rlMV4sU0JSfgrwf
fqxihhxzx4VcTCXKygGIwqABK0bbtfWb7UeIIc0wO/UOqh0veTHMAc7ZFxfQemupkYwsHJYSRq9n
7rX/jRZ3G5oUWdk68f84EgVXJ7WFuQQnONBG5dRwwtEAp5sWCpigQr2t9FI2b6RnFRqREzb/YOvj
hYoYEVOskdkf1nJ14Rrc+xmHLIS6mtMJqhWHyJwHb2PoHhM4RXvvlhb/uFrBq2qZMdJNMkIg1dQr
05PAarYuC26bmr+t5vpy/Y2UM2fWeIHuiXLR78EB6maVwdD8CfVal90ZUC1YdSMLZSxECQrnkDm2
nCp/HYUWR6HeB3KoZo7MIRRQOrwT5TmWrK7YtJg4DhQ7nIqzN51x7PxDfkKPxhunm5P3b53Noq/o
1dCHzeCQH1jkti8ZUqsrXJDzL6B2JOvAQm1R/RaG8QAYShIP16ECjj1cvyCVcxWTXNsBdnp/Oc9I
EbfPJEUq9HL3rnMmY9N7dJgQmJGGV4lSVhS0onIHOwbhlOnVh40W0NoT+PqaxwiF8ZgvzwV6Ctrf
tpCuSuZoaZXHozDDN+eOO9zn2ebt5cXNFK+tpbocLpkWy46VeLWTEs/ztzcVW83/FBKL15ip8BnP
pAl4cA23TvDdlyOX+BnHpSOaiMEvfS4TSaugyBzUsltaDvYsZEWNmMfVdr94h/VRU4ths/Sw04YA
vU0qxi/H5U8/U2V4nheX4YuPYhcOLKbYeAu8RsgYR1PWmZJxLwvFa8BLL5Nw9CIiVKtsT9TxLHFv
nCRcZhO0DNrNDKaGohrROngVPd/01aMHXRVHIg1XAAmoFAG0Br2Ir5k285oKUPfkTws8OABZ9rf/
zEMXcxUqHbd6rHGgxtPi9KnVWlP6OAScb2r8jgJy5XSd6O5VNUCnMSZ7TBRAX9tn2hS/rd9/JRFW
QywIzfEh+PFTqRqijKPeX6ivcQuwDYw7qS94OSlKOjrXpK85UXyc14qrh7j8USC/rroSTMURRVox
U96Nc6/5rTdzrzHMVBaFQZW+UznIBAUaVFA2EWpjHyGW9FIo2G8oo2vDkIx81CJHsewbrmtcOizQ
fl5chcUMxG2XKwqyXUIbQ4m6JcXlzBT9pvBhg3UK9nDmkxdKVgvyYRK9lA0PZEZCpi1NdD8MtWPG
q76pRRIfNvoOV+ukiLT0pkgd56Yp8NxRWaBmt8PSdKamnBsCnjVUUMMbefeeRPPxH1vKHm3qHo+T
2oDShgi3gLgnjCiLoSduzozytS8+8qZsHCYZXRHPbHTxmanRIkcxb/0uWlHqIc3U5C9eajuOJJQl
g76OSNgNtrTyv7ZbGsuuugvYORbVcOYMP60Ctgb1iny+h20E0lqGcTjYw2VtVJkjxWkiAPIDGe+Y
6HVHRMYKMqPUTOZQBmiANvRxWL22TjDJtZUvNeHw5jwdgAgbuen0BOa1WjOUG7JrNo4V/IlhxNrQ
IfQJj/H6Ctmi4lMKCNGU1UyRnWsAFziZf4U25TGT5gutdcZc89EE43yGiYRZVnzSN90k3pOAZe/X
RJ8Ho112pfZkFQ/yMPld7534InbjldJUx2dSng4cqa3hJeD8fWRqc+ShAOjVZL02fCc+pZdiQkmu
NOJvDDKcqzZMoAABPKTZ50ixuG5BesBJ2VNZHxy56KaGP4/G/7HDNETBNtFna4XxNfQ1s0g5+j74
aloneIt0P7HgdDNLUyISxxI3CX1n6CkkPuxFewj92p6n94iVeWy3fOt37pifU6SfUGzD7gCQ2n0m
ph4wiw4gntaR0p9MZbcakbsH27mFhhppZQduA/Xx1XhvLtckDccIDYXxgF123OsqVejDzFnFH1WI
1b1IwOAKV0gr4IIW5Hv36IShbU+AZZBffvvZPJ1MK3ejJcm+NN/Sr9Ul0Uz+coMAogq1ynCDMKt6
G8YqoXyHV3jr6GqnK3IINCy+17DiqGmMdrwI/5BUXUCo2gXzCz9WMjUuqpWgFmQ77cqQArFoozXC
eGNNnv4UQRPqFUa/bwQynpgMXcxOiOJ3YS0jCno33aY4K1hmBlLoA6fHnQd5XQ2FeYsrgTSCQwzA
dzYw9OFX5Dp3NMsTAOkWF3njp4nwHLCFzVy4I0+inNl/OQaeae8hSfC2eUsQi2pyFzYAvwO1AEwm
9gRQk6OPG2R+W8k1JXCLx4SlnsPgd6DUZIBM4zIE8f1nFP2xf7lidQB4q95aVp6F3m5T1df8UPEB
wg2ht9A7ZQnX/2yzUgyXfSL7ZOL+jiPHJjUvyWlRtuRHeYrQXubQTm4OFzVKlJ4etwQjZTwv81M4
KdBTcmByq6P9IQmq4zS2obVu9IE0gDA7AuWgC85MXMsHYUPn3b9BBYjWmYO29WQVcJjp9j3D4PIf
n/chVBjtseLrx5W4q4wBZJtwChjRgWtwmLvv1fBW+V5avMKZhKY/cUEf7lG+PwCvi4Zz7rPc69aQ
EW+k96vS7JzAQQ/hkc6F7zm7QY5aMBVJVJO9sw5H2+lwBu/CFCaIBp29mv/bbFL4fpFL6oVTFI0T
5r1gWft9Cn0Fs8peqfLKcmnpdYriiUp7LVe19Rnqk8uAP5nmt4ZOrc/CN3kpFNY5sjfRUp9WfBa1
g6iP/sBBvGew176/JXfoc2oCLF7X2uVioLcswty197YN6UkVoLgUXszEaPjtMqwXEk4sZSkD3A0N
XQRzF7OLPgInX8VKylHdujf71PJB2cp37jurpQMpkgi5jlR9Y1vWXx9xjlNgJSywqHoZHSsG88DC
70FavFhJv2E2Sq0pv/3aKMHnfVNjj+4Bxc8UUeCM0aqaeQkw65jowDRTIQ7lo6ZgnUUeqZP1MxYj
LQP566LDbxDUV4dAa0xSL5JwvR8KyB56SoNvs/+A5BNkOi+W8hQuscqsYkgVqWqaHBuwLKt+Y849
KhMYjGTjEn2mHTViN7Vz7j1hGf4YF1/qmOXCpQGTLGMsDQqhHbvVXsiZby1s+VzueH7IsjDK2aG9
IuGyVYpynpbzOAT9ciIbQOPOCdHQmIbzsPisNMJ8GDgvPyTl2PPL4XAPhqbKViIZEt2V+hIOWq7e
vOLB0bBoSAh1pmGWFZhAi4jezXQPPo7zUwnR/Ffpp3gVmO7GRWGCXP7+/okS1tmu+8zSha5xbzws
3EQ7IJDl6ydZUHq6i7IKdbITAAepEpZGz49/yay6h1SGy6TObOTARIdGPTheateQ+DP58XOwOlIv
vTZ8U2IlX2+ElRHSsZ3eqPmH+e/JXpYIEADICAnteLJMNhJtnWVUkh20oJGEmIz01LQNN1bHncK4
LDhtWvSxGKLa3vskLunTS1fpkV0Osh+uzsQDc2Ka7DnYehAhKJJ+ysbktDv6phwyE0zgkyAhJIF6
0qjJ1lZa120NfnxnZEYQuZrpZaN6hcNlfjt6CVGc1XIG+spAUCejzP/sjw6fzr1N+I26FDL+z/BT
w3iAXjLK9rXhcr6uBReOTqsdYVJ7lniXWxn9YU8/Nne8yi1gEQYTke/CUkzktRffdcATslJbKnK/
nMhm2wLaYLurm963byCmQJovV/ABP9pfF57UdSTnCHqUV7MhqwA/9axwi/LP0v1CfntGzvXJBdO+
hk0eImtS3IyytxzGKS/MupT0ZBOhdvarsAzwUy2M5d9tinspPT/yOOYtLR9ilRrxztOhtD/TYpK/
acjsxf5SYsmGBJD6PjQ3PlINStAMH3t0yVuvOqeVXGpb916vgNrGWC+Fr4PoLGDwbTUk/JQuwjop
Jk5TX+gv7TDI1iMzUS815kYQbLfHvA88T3b/RwXSM/La+lOuUFe/7I6UeVYnvF+IC0nix+xy0kRg
HwmZk7zu7t1PMLaiGE5Q1X+X7Vghld4wvXhEbZ8NLeYFmCw15Mjy31FJ3tkiPzOBCpr/wFqJae61
bgekUv6ApRcaKRmTyrQWKSyphHwzFuTSQkyBzjsgQLblHQDPsk64/rDGiG9hSsaOXrJxNtG8x/7G
HCcYiwadJe16vIl5O9NB08Utubi1bcM73A+kvO+X5Q22TMU9v4gKD8ombTtdEjJUMv5QblaDWj8O
KVsqT9002slhyPduDmpD3TMu3c1aVZq4S9rQUlxcAAQrtwN7X5zVwbZmWZSdGnt4yG2UaTIfi1H+
h1YC617zg2Dx6YZsHNcjBaz0gDLrpBVu6UWnsmvUMXSVNbThymX/0LFZYuowplQWjWOw9CZHgN/c
pTeJeALk5eAbyn/5j4i2fjuxpY3DMLGwuNDhAMCFwQLuWR+9Tgywu25GhGVna+xI0ccqChCEhG6w
/1iJAo+2th6ZiUvlxLmqwyI7XhoaaHHiUTD3lid+km+CODd0IOGuxnzoiV77DCoi4WevY84Re4Ji
iQk8hcqPegHUm5yLx2qrI3kGevNUxoebUyewm5tRICbbEGMSx5igncwMBiJuYxaX2ZzKTm6V4ETP
n75HaFQYoi00fyFYrrQl9R54QetwxJ6vJ737sITf9qAFyISSqCIN7SGRo3aDiJepcaDxzJlCqGcl
srT5br+R/Gz2Dks95VK33ziLbRd6WpSFTKWvgOWNWV8rgHFU2OpgA5JqEtnwwcEgypKt2lkooZ3W
8GIPZB3tfCvk+UCos+/ewtMKcvBJq+iFgQktdV7R6eFmLLPsurLxThqzK6meZNZkXoDaXjHLyOzi
qfH1fr0fhK0nv3Ey7Efxwl9wLpn8CPhIc05uHkJ/t7qgWfZKhfuaz8jY0C+nxxbgRbL+g9Je4bCF
GkcZWmephGGjP1jmV/rt+ViL5mLqQEx3IWXsEn1hqvINpMvhDG2PgCSw1e9jB2n1wPxSbhyG0yMw
M/Pl1isk7yF9+JG1MKaab+jIK1GBfmTAYd81S50h5VlNf/z+xFkrD+NxxMYmObOXUTxMuUmTGYjj
dpK6ZczE4Ysx2cJtGxZnQ3m+Q9ims5b0Sd9Lc9dG0zwPkS0gER2JfvYNUP9W5JX8Im2YV6xChdE5
x0kg6+ornL4cdtwL6VeQSJGK3gB0n+kkp7GHnF/ljSZ5yYQIUG8/ivJ3nMgjkTI3DfapsVryw2Yl
XtscW9b6Ck7Ywc8iqXASIvQSo8q/J8kwZ15l4T89cwACbH5zvrSaiOdwXUagy5Vc7D0tx6dYW4EN
O+hKCO46XGLHrPwBWZYpJBv4yA5fJzUY2fGEnKBll0G42cyQIM2rjCFX3MxrYh9mWKBKwHqd4C22
eGVkb8QTS9YsNd4TAYMsabvK2eymSL9J02rkuy+wocPOLKre3t9emEfucIJB9GViRs4bOSDftuCG
ma5ukj6k974xB8c659EcW5W0xQjys/EkLALKctJnakYScoHqnPuarJZQQXJlDDpuzDbq4fp8psqD
uE9EK0B6Ch6yE7IadEXSBbXWj+EdFyTS+XVn8wLyJ0IYNcyG7xrgpWi9/A97xw0ji5BIq3vzdjEr
d4SzMQ9EYUCEXgj6RF84qfFLtHE6uUqPLIJ8XS2KzOEtl1ZqAhuf87LGbdZJfxQTQl8Wtw31s16b
Fee77oiyde8HdaZPVmzxLKiPVJBh1SvqxFUofLMj2KZeOAb7LJhn+o17UYbuER2xdH2GISOgdzdm
MPktzGaGzuVWpGXtTFXIk8qamPuM6hpb1I5UfCFy6tMQflEvRds0ZAJSS2CD9qTPAheY2TZN4+33
5y0oYvohM724LyhWaInchndNKmLc7xRqsi7rWW9wWuNswAtVLbSrDxPWaP/dWE+/5h/yXVHbNyO9
IZZKe09jcJt3Roz8wiwNcFB/EdaAjNN3Bk03J/ToJ+knCIeFtfeerMb/OCdqX9dqEl00VPt491GS
0tLhQCwNibqTXyWT6dkh7dmS3y+usTv8aiGM9Ft0l/XRpdYsXGyHF2HkC/gF8b4cEYZutYcNQNr2
drD+n7NPDF6ZdW2HTdjiMRHwbPXPOaNVEzQ+tm7n7PJPUxYeuXxYEJnH2vG2pY+bR3QlPT8ZqNe/
Tu59eHvvQa8GThD2fWykFK3WF0DFNdGGBJsmRQqiimfGY/P9cphaUuH+UkrV/1k08t13NUZudcRP
ETmhkpj7NYoe2jZhRpP5sbCF4F+2NWjtIcj1/JoCG/hVVO7Ep0HyKI1h9xPgZ1FpV9tb36XiSBih
47mWoEPKgjAc8aGS+XsK+8GxAHYJIuhmzvZO65gA3WEYdH62y6blrPxpyXlNuAe7nN4bV7XSS+WQ
02mFrDQXFUZgbgxL59eFv7fom3XN+mXnz0Xlf51q7Rdv/c5nfD73OYlgECRG4aDlTMkNlmXdwqd/
ylAm9Udx+EUXGQoK3C0wJLmABPkzVXWtf988ain63R3AT7DrIYZhb2IbEU5Eo9ToT5rY8AbepIgk
Oh3bPa3q1Lvaa1IJi/oCan+6VmVE36cHdjTAiyGg26v9YI0O1bGhfYtBTnjjP9Pg9g2Irg3l3maL
AngYvSxeHB5y9ojTg9q3VW86AaxFvVzBnT0LUH5lAabQS0QcGT4OyD98xx1tU8Faf2en+TqjuGYg
e3ny4LP2GMk9O4THxLPUjF+SNZEqqBGgGjYqwoVwJeoOxqaramegidNkE819sjTZczxyWZBjvkit
whMoI7injkOgzHchFY1f8zzYs9vLx47/zJsbx0GOFpgw5XxD57+cW7zlGrIlf+qb8PwGiEntOamG
ebm2AGNi1qf8CKsgzDumzT/SzYJT8rET14iw9glPNZgjMTU1MepmnGlJjdlU63pbDclg8yQ3cRgQ
32MS43wFx+xwgpU4do8paSon/qwvPjB9p0ldCIgqL1cKDB6MYjpD63kHjf028DKbo+UO29w66KuH
FFvOKZV6Hde4ttBZI5z70fU6tU0FUsSJewChso65K64n2L0xw5sRBSLYzkfRNtlkhwz9AohLP8k8
/94SriDRq0YEjwEbfJOF/0OKuhNsP2OyiXEL8LK8ynzdd1s2Xo5rClHhS3aopZQYHtvk5qa6/byb
ty3Xl/0dAkTf887sqvQ+XORdLCAXS/UcR+v9I9nli2qgg4RD4gdb646Zh74IJRBjPRZ76yIrcpXF
TyOOp+4KjqPCkFfqYHNt4smr3Hkc3HrSuBCFtvuj0w4vQRdoB1gjuJ5XGpkR0qpJm2DfJTEOUiId
7IaBpGekpbNyMlG/x7ikorJupPz1V42/Sf9u3MG+NlCp18T0hpzKr3YnfmCy9jgu08WhW0JmEJ65
mQIPleffRS73g8Ap34xFvaZg3Ee+m3hslioRZndKKKl9l73zFivVwK3qQwNuMByEtltWMHbfRwjE
ZF/SYENvbAZTlLOPwgA36AcGAfgl5HsC+92XnhZV8KtCmImb9xHNVtx2mLYA4fZ6BsqkKead0vKI
YEjtJ0mXvfDiwgNCnBd+3GtcLqvj+mSolJ6bxM/yWsZozhBNT7/XMupRmDib8dMy9ovjpPg+VrMJ
PlYReq4+O2Io0Q/wW25aaCWwqj0EADwfTLge97iS0keN03OesWwAWrzV7QHGPHgPq/msZkUQ2U6f
Bi3QFC5FB9pgj4wDzR95WrxljErOyUvysyNFgwdpgx/TVw0AkEkporPPlXqiCztMn5zydVk8zzjg
9kKPYPySw2+z2veN3YCiDn0is0Qal+xsRRHD47GLtX8XHYsBNxss2rcl+nw8WWHnrFIGhTvmSswa
Wri2YSQHMreRE9QRw6LVUXnhZM84/CD5aLmvUPU8DwCeeM5tBU3T+MWooDdjOI/+lJZ0ezP6fjZ3
nPlT8+Hs6P+hBJsJ9FktVtuKxxpnE6GhsMaCmzj58xC2R8/9Fy4wuAfJzm0gvYI4zQGMDa68jgpj
NrqkgW8PJiCLTMdU0iui+YiBmSMVuQDrc8v872qGFBY3v/JRAbDUboqE7YuZHT5MG3CBYxeo5igt
z/mOIUfqEitWIVd1QE455PbhcJQS4JKZs93if21E6l/MGUzJKFXpLMtLfkG733KFhD+ieoNiXUev
fK1ql44PDuCPASs4BVNZw2v+3+gtk9aowai6JuLWST26PDIygwZyj9sgP3yGn10L34kEBlxLBY5f
++G4Mjqh7uPRzHPg7sQTw2/lD4q5uf3DKc2ZCdKYtpyUW9EIt4WAAYXPrzsN+LXK55qjtdWJgsHu
iqzvgXowlTnQLZlHdn6i2FAYVk3DqK00bYMsKr3Vlxys0sPbyqCOmCI9g5MkmApFiMWwgInsqKnF
GKjXk+h4WahslDsPDSjgnEcHFl5tclAkwvn0dc9mMG3IEJS723XcbZA4YQhzE1aKv7TOHMAr7qFp
gRzg+nC5VfhouAP5wBFDquJyWH8t6EiDSYxzI0HeoxoXa7/17Zdm+Qmf03QUZDgwFfUWnTARQQKA
yJs2NzK2LRL038xpDWLCp/frQQAmG7LejBuvzJJMcU4kyKLZzQr+riUcporqh1AcPjajQp9QZXd4
1ZFSc+FBMxN9t5+0o+x+WkY86neDDZKwWpGFTGfbl5/cn43M8vY+rD5tYvmZz8bHC526g3w8oehv
GdzaxaLiS1WjJbKf4DJQtwEawyTxkIv0ibDb6AZThevUvdX0WDTLu5RZuiw5mLiH46MKfnEU3toQ
jcYvZzsvpdB+vegZNZX5xAVhV1e7uCd20AhMqy3D4iiTe3CLH2ebDeH2Jg5SRA1zM0RGTehbHixa
fdDrtpQoCZmS6wLE/beMA0jNOFIUsuHvEUdq2sWzFdI2ecCEI6ninHWUQ9xRWEwMzexO7PrSzmSs
SZ0nt1ks1b5d5/JtSpAaPRHElkxabN3oOpJpiajddauwJDHRjGX2XFMJhovhCvboqLLzwuEvbwXN
0NrPDKef4NILZZKZSkY8IPR0muJMWzfVoNK8CLs/d3T8FGSbW978UB1jnDk31tV4YO8cl9cur+Ia
NM0mnOhkIhGbVJLzDux/xRsY/8vE9n3s/i5ek5yDinDSfpMvC9+7zB6qggnfBQwZhTSiF4cf+fTy
BIwswRheDlN6jPS5Q2lIc68o/ur2tu9GRBCi7YAx2xVsFBs8z0yiwtJt9nqLFQ9oHy3+Kr9u+EQ3
csHESCyCJyZUg/Elr/dROyCzHXaBrDBainmtV5dKAPGNcKa6xytHpTFBDEq+he+ZnAYhYJcbWmRj
7lqfD/VrnGIcOBxhYuudInEPuUvKl3ubsdTfcjjyNDTfp7GY54UPufP+mKF+U/UFIRE7fgK7BbrU
t2cFjiCWHzxGIhwtmCtiFUtZxCpWMtRrHUvhD/qLZ3xvZ1zd7f9fbdJ6gQrNxOfquPnrRO80h/Wm
PqOewrsg4z4wYVuAZ32wu6QMZJpSK90gDd4taLLqD1z5Gl4Ger02HvcyvbO7mNkTI/g+KUayMfh/
iI2r9gmTKsO+VEIKqPw56cN2BNBZrrb59jkNM3kBN+HINDuF51JTw+eFq7q8C2ieDBmaZnuxsrX3
7fAhRFiIini6D5aXQq+KL+YI5w0ILpS3WoYfq+S29j2pD/N7fEdXgNn3wMJ0MJ5giQ6FbjgPiCdw
U6ND2t+RYL7OkbrqgJRzdpWL4+hZWIIJdLL1y0ebu0Q42IyijrIrnxyYxhAbM7wp3wwizKiu+muU
daXHEUpWGkfL47e4vSkB5v/7BEit3jIgnhI2DQZmcCRuHMFndOC8KmHDOj0t+ZIm1esTs6KZhk0l
AoiIgbuxRzXJX4Q19cijX9nz8wPyhsByIj/3h5ArIYMQwg8f5kfRcV7bys+xM4AGN90sHISCql01
wd+pp8zbGlwYCCh7E0biaCW8C3zoTAZbDBmrHW/y0DITnd/DlNeswKxIRE9ydKwGqLxVbJuXU4UF
ldeU3seWyIJtJEw5qjA2Dk1LI9ZJ8+KF2fnNSyFXf2v19onl6DdkHJf8QQBp8QlBQSwkcOEJsuMP
DJvdKdYXWHu8oqgqzC5dn22y5ZyBoCjVdBxp2ArTRAjl3oUWGZ7UI/qOENTadkNjjj8a3CxNxamz
tJejqZCK4PHsPzyF6fWwDEsINhVGTF8bXChb8mA7i8Vg90qdrYKVbsK1vnPNKjuShF5LFtQrrqyE
VJaiUs4Zb3VNCzQSrcLA0+N5dQcPEVz3wu+iU0t8hLsRuIhv0yVdMbf2pDcXosR5qVYpKTZiABsk
o06HxA5dDgQAZi2aQXQQIDcpfub8DGcasobieCGkxcWotDKkM/0nk720UdqgJXOvr/cIWvc+HC8q
XUI+8oAQhD9Dy3YfhH6G3noH0SmOo/UAOFo/QK1AJgj0dRDKxOXOo1KEKzSmO9luBJ/jgXcczvld
qTVQLz8tnkRu4mbbCRISJbJQFr2qgOmT998gmEQm49OQk3NSE21UPs/OUu+M9Kvkc3B8iHOEd5dZ
TSdtIo/F6LCAhkwAibMOMHnstba422DNuBgJg1wyHZwtUwCR/j59g/Kh7KtUxtwLkZOiqKQXMi+I
t+nBwfUTY7XgTOnhpEn5uM4moMuL9GNMHIJb6FEZi3zJ7KOLCJL2Tvdu2buIRjBtA+L0or390ZFd
2nDVb7kVg/kOnJwVJ76di9P8k8/3/30aYiGoTH/1+qkZTg0rwS0Xr8zz5W9DZGYDg8WdcnGm4TJ1
wgooK898p8rI4bAzEcJvXlLds75pEGTymPT6R57gW6nDn2+eg7Nr3PVFxuo0e1uFMugLmQn2qABb
Ym3K+Wp1eOOWTTDmpNm/eAdh9KQ+EFJqQu/k+gpRKGipKngm0UoThxmY49bUcpezjU8vnB3/cZml
3KlRo9MKOstbJKXnek4CDckyqFDSyN8wzoczIT4Stx7O0aRL8i3P3EeNSJdnfGUCOXhaAATXJK5V
vh8gFAm4BoiPg4mHklvBu9Ul1/awxEwoVLIL+qtwe2ymNa2ePzdrAjNJgknwYIvJuA+qNCHD0wLi
7wwEXsEpTDOrpUY82obl+4TMQ7mU5II1/Zi+Gyh9knJkswaQkOL695hNf5vXsSMuRLdFCMI3C2GR
T0tok3S0aPuDjOmiL1zv2dQMb2UB8RERoufT+OSEQgl5vRZkWGDODwYjg8vsog8PgEp7YxUTiOOz
Z9/1nYsoBWyx/K8jmtQ8HGUJmdM91Wi6weCAKbyU9mG032nSqCV0ZYrvWw4kSTtEjhV3IGcURK6R
LjIJ5IMnsLBK4GvYDcamyG7M96tpYjd+zaEJZ2Dx05O7ZUoAK42nLcll8fRamXeHaT1ONUb4nlWB
+IoHQpiVRBYPu98l3u8Rt6HS3wvf4eDIZ4Hgo1YrN9uSi6L5NM+oaCFs/hRG0ZZUU2eYo6N7z+IN
5ODhl6QG8tgIE5zLjAZR3bbWQIpZQEXmYGdln9QkFteaUS7mribH4wwCS9GhzvAcCuaGLdapKuId
MxXmrXK5ETWAAgFUISHwmwNe1YELALA74iG3KrNszq3PgCO2Ci1qILolTiiadWoDsQTtQ+MGFWhS
PeZ1xE2h/NsRPsctFURMECrdqWfP/UqZaHvgeI50QsdD9KR0pn/vPhyTNcUjtNTIBdhJFDp9O5EZ
LvEnMhHU9NzFpRtMEYZEMdJ4TM9LjOfTY/YI4m9Z2UauDQO0i/QoDCJ+4HLdf6B43EvLQ6NfTq01
7NxCHJsleWiQWTIau84iU+AxCUehfwP0H+l9mVUZwlt0TdNsPDsP+jw2Ds+U/AmLxu80zmD+dRfV
MSiXR/Da4y5zbOm9PmodhDnUmy+HrLqgIKkhXy5fCc7rn6IJL8buDdmHjcstiJuHd7/ZIe2qILY8
64nbB4RqGKYuHD+Ioj/I247Vl2xuq0MUFyU39iqgFPMbTscEdUBL29WCECVkNzp25hQqELCBOWLV
MevkFRjlxEHgImSoO+KybdMS0A0TemjXCgn9ZBaAFBK3Uzl0MCFm4+BHDAkJQBdLCsN5X2bqf7sV
+4fU8lD5r8NesmBratkVykcNieCKm1v8oL1nBx04GOhZXVdLQjlfMaYwPXUp/Ux3yRCtjb5982yK
uX+1/S0xk2SWY/84iOgcwZKnxK/uGMAergkAfc94dCzM1cIZLBq0vqjPC4bf2L4VLzCjq42eFNgo
v2I3mmPCtc9JW40a/HiyyRZPF+0+1sZLmVxK0LSfk5juZoJWSa8X5y5aU298mXgxceLlGF+TRwqj
T80nhXiH8zcQlP/9saYeXxDY7U+1Kyt5bd28Uzl4g588B8OmraVRuz1xQbmZUhFFfesTNgSKmiHF
V25TR7MhB6EOUJFv1lh6Ngt3nOCi4IbgFoD0ZJHkafG8EWM2TqHI0XqQqpTvCumtxzmea6rg30Hl
UFWw8D481Z8d2xxejaUikLK6eJcKvGR0OCOb8DXYzCy4DLR90KmjPlwYcrcavS6j7vToNSzs+Bnf
qUZHGnyJ2QyC9iluNZZ0IFlWa1zV/TJnXEpaPQ3EsSTt55JOCS6jT45kxUTPB+VuRmz5MbjTVU57
b0AojSZDSUAKhuIX4Pm8A0ti38/DHtQkyvoVs6wnh2fODrpv15ooFlaP2xQ+xTcOJ2ptX4NqRcKu
3+R1ff/je9c+0GKAFgsUur78lFIu8pfraXm+zH3ihOZPfG4R7XxJcbK2gMJVp/1nl3IVuqmUVLs4
kFVJhrUlpcHVKXsZPhpnXEH/MQGaT2lv9qLDL80ene1x+WCMo6VWX+wJThhcqe5GYGbbwxANLO+u
rUOWF8ZpGGQKee7pndhjCXNyi/OQ4pAQ2NdiEp4LWEKfnjBbVTQii0Hfag1dTCgAUEvjnCTz+IDU
CU2lGgEqz2xSzcxNLHK8MvvdA7IPJfrANYxFecjbKZ90EKlhNEOuLe26CeHpLVlMFXjV8NATc3un
kiUvMSGAGEuP2+NJjpfOxFTjIENRyctS5E2va5AZkT8E98ISjHKEAtjVOpKySDBtcbKl3VG1rmtu
AfqXauFAyGmi0krieigmUNQL8T+C7faX2zhfhftkK+Wcrp8ZsZfm6qW99T7lUd5xUAn3bIsIlXdM
wl1HF94tYAuNAEHxMqRn1kKE36GL6hH2+fvDxXZI5NVuF/qVvIgtZgrQF0ZYx3Nda+5RROAfG8Ji
OcIHKRMkbz7wuNika2vBpTDp4kPLuQOqVVwqCtvunaCtN4UgvGaJMtBfJX8wW6jNc5IH0l9AgXOL
NRseBPTdazkUhwKTh0U44CDJKiMSCp07Q7tvYXz5xyAdWowsUljHpSh1D+q0JOPy+zpSsyQQbWT1
We5if9TZ4UNNvOki8eUKPP8un+nU3lN0uR8f3L/KX7Th/KiEh7V95qn46I7R/cD6IxFAj6poDGhE
5WSTlIExDLeP04SFXfm5NjEgTFcq6gnI/9ASvrSkmmO4TFReP9k4JNj79649JJlgudxbPA8LcpcT
KdIxwYcLV0HlHcLwxy4zzu3JxYJfmUh77p3/ncDd6HvZjJVLWRe2kw/6ohp+Q8Vm3y6r1zRkcgeq
pFwdlYVizcD71aNFAJ3iW/E6LSuGXof8no0ztpL4ys8CBbWLEe0qKjDazuCSjWuxatp76nYgBEFM
5eK2iZK00gX1oCralN8JYZlWFnuRmKQ6zBnY0keIBLC0kBbW+gcBX727cjghTdedLR1k9fFM9c3o
sOWKL60bu8gJkPBB/dQUluEMfuRHfCdMXoMMsei1uY83LFrDMLF1o/KsgOqv1PbOuDaq91GEY8o2
z23mR5WKkxOY750yzauighCMYuBwxqC+3BUNrR89Rc6hRxQX68MiVJkNwlhGTE8crX1x0Fnc6xHH
pdvWbLnaAe8OCBijevSZz+PvwMGw3WxM9Ft/XDN6rW9ay/UxRlB3eoYGtiWBrRR4LSD0IpeGJGKg
QPX8SpSjXyvqvTVEWt+dRtjc4fAu+EoDJGhsTVIn2Q2egyC2gFPw41jARNCQaADgXwyQr6SMkqUQ
9qnvTg1VvtppAZevbX11GKj+Kh+NlGUiSQYqwDqrYV2cP93FY7Mp2AxFfZT9UoA23Kn7NzRS3THP
UXWaA1JdAsi+QfwAfLwTLoSQdll5orYppDbEpP84lFgjw96/fceRGoLsVJAZABehURpeRznHHUy5
1x5br60LqHEBDs5w15JdoDdHbOAcAYGWl+GArWomKMJaz2VL06nN/5MzYZywKdYIB3IqzVhFhU/d
BVtYIW2OS27dYpz1mDPyrHVQnR2eS++o9VSDhIX1s2Pm8lgCGjxYaniX/bZ474QFiXRkUlZ1kWaz
Ljp2g+OOzvrcF+dAZ3fIPSQcrS+F72vciOKaK1ZKA3jS8kACHk1A0SGLZtGUcD/8os4Wt/7Yvui8
xTK8w73w7CVDZAHqTyTNBk7wuJLezdAK/HBr8ovXRYZK25fppYIA7RGZLjMk1AOuxt/I1ZsZofJA
nIBIIL7B4+ohexKFHXRbOUiWs+4T3Cds/b7ZeXKvXMghn4DvABLTX0gphz394Q532lTKsvmrbR/p
wxtypy+R4gCjt+ZyKUncncpShxj1oNJP2kZ7Lk6YQjk+Wf13CwNtyyMPDY78sVcXSzgY+sYl8fRm
Ju3xc/Fa3HLcl1FgCilA8EBFftvSySDHWR5y6i2ntmexg3eBpTHdenDq0aNCs/5v3A/NWQrBKXkk
g1RFAQlVyYBlA7l/curCfyqgn1hx/brKI2dRdUfUE0yZ9h2FWYhyKzqy9t4+uLrZiklVc6texDW/
QnXogdI2XDYFs6j5cX3Sc8PfdK8KGc7/Wpn0dhZ1x4ee9Qo/jglPzlcrqGff0INgNuccQhoixy59
GX2nevGFINT4zPLjuxm2IbR3Xs/jEOCykBoHKGla9Ej1VcDkqmw3ZGdGP9DgoQNxEC+1gj1rcTBJ
7KlJ/OwSKSelsBIcfdaXoOmd3yjXsejCiZPT74CFmKAVyQqB16lS5zsqEjyz9yD0xHqBdJIQh38J
8DYV7z/WcJubU9xv2kbrNUo3dSnumdyONQFWTMfjKDQOznYExusymoaNDEwogpIy06YvCE2tJBM6
3t8/2JyYlXO+X6NXEpjd/7c2esI5VsOaaApS8TXWrUqDcQa+TsBsW8EmRX2JTx4to5/ErOQ6GJml
xNXg76oi/T38n5dhb/v5MUniKzmg/Z9PuEZUgBA4O1IwzFf7NTIvAPEvpsCjiq9DYTqTueZcjMV1
LB4hX6rcLOKK+92U/7HTnR+DfWN8m8Qw3pirp7apnvDPpCRZij12F2gKjKJJ8H4zx9RXW7T8/HVL
fXpFTbWtiwZPCosYsaRxFXvfXg82ttaR43mJVRjUsHAd+rolMEjvPRWECYKk71B10BuEy+d+2Xr5
j1KA3Rv+V0L0oH+y5HsDIS3Nqfv1+qmvR1SE0iIM7auEiPup+Q+sKux8q6RgFDzaBhDlXJ+Wgb13
MNsQs/0ztXVOdDQMEwzlArU61k8k5nXASC4sjb2E4WbljKTsx8x2451UeU5CmFBrbT1fKT+gYnN4
DKbaa0Z+PiSOZLjzqA1qz0vaMgiRPyQNadIyMbowVXsVAh0bjmUq5agZS0a/xQSKyvcY8yKltqBe
zeChZM2LAqNmIHNobF6D/Sdc3+4uJVKFrD0blbIYcq00gdZeiPmO/PIZpnO9AB8Fk2iOd42J7KiX
jvgMzDrOmP1DYTSc2a/pXvvSQZalfT72DbSM+R5CjQ5/CZEMhg0kBhbG1OI09eY398K/sRFQxp6M
cnzzZjjQkwRAIo6pi8nda1j2M32BmXx4ElKSUrFZTBAr+m9jjp3UAsi5nauL/E6V7lcwTovcxcli
41hx9FszyBjFuNXpC9fIiYk2BKnmKK8oDIs2flnYkT44BUa1Ih9RKeO24qt/lra6DsLMUGRCxgRq
86DaUMEf8vzFe8/oxq0joWWlBWA9pnF2UG3YD3mCJVzVGcwkghPj3teWadF1Kfg5TZ0UXh7qsJw7
bqXP9W4PUDczLECAF1we0zqHa5SpQj3HGGEsqTkLCjOKakWPCpcjX7lD6JpQxlpe5TnM9PBLk8eV
QWHQ6BxSQlfXlLpL6rs09HCUVoqzafVbZQh+yG2kdtEzRgnXZTskSO6LzMdZ/M6/VgC1Imi9P7Gl
BeOPRC5VumX6VW81eDo4MypW2lG1/nZdIHiafDzreZAPWzBp7hE8mdB4fuhXoOj4SaBtJyPSQgoq
omJkQNVGcJhdhbmZnavtVyLK2JO5wUmBP6D3T9/93LFv1TJEgSbK2nwXjs6BfdwtFAyLAYSZ4G0y
CzejBaQQxq7LnKYlBuwBrjwjXvsJDt2wCVuG0WyFgiGFtcVewDEVAP8Jd3DUBGvv6SuHKQK6SuuC
ZFWyGC4+3DIEqG3JmESE+wuvURJvGHBgLHrCr+paur+B4MTUMLJ076Y/4MjvabFwcEgu9trzYczT
fiHFqTenzSMg9Z/2hHGfVu+XPocb1KN4YHQ4FTC9rdkajRZdo5+Yt2Lqz6vCZqmkTRg7rjjCZ25q
BS5cy6agsIMkCSPUP9/oEDGutT81V4IOZp+58B71aD2dGfAI3a7/tSrctXGHjVJp1BCGKkMnaAiT
3lcphxYhd2IvnGQRAKeH+YOJcXYX2qQBxN9CdAL0wUexUAkh8xkCFp1PWA9mUiVzDSZu1PpYCg2g
OG7vKWQqMT9BDCF3R2SS8txdJs/jLzmIGBJcLS7PbFuj8ZJN9v5DZM5g6/X2N2FWdVcj1CGLysDL
HajLDngMgY6cffiULpNwgNqwBqiDHF+std2SvHYj3/1AymVagYCi9SliYqszAey0hsSJ00IlRzJt
WbHhBK2fbpXCj955yUyV1iisP9aT25RFqmJ1dx1qXu/b4VFl5xSIJch4m3FTAmidVamSTr/y4icx
VfM0bFlWCd9d5xNr9NJ4kOdIDg7//NdVlMH9UUGUzkBTtUAM8tdKPUVUuO3VSIw24sTFLkS0pVvR
r6XVL4ZzTrMKOTGnECi7VFZEulSemcWiO5FdaNU0xaUWS+WH+QJvOFF71IxFz3hvqNCKUeUQ2FOC
r+pCWqAbfn23y59XnlHetlAHoRenlr0QyR97y70J66Y1cJKmWqof6JbvbkYlkm2SsaK7xkiqLhgR
uqfdfgF5aRnEW66Bb9tDM+MjBJOvQujjiFPt4fZOROnpnoee/PzQMULKaFpqRAbIMiIRVPmoZHLE
+oJjBchR7w/6WFoHHHS1YeY0nD8XwZ2Xgqm/KRuIbuwtsSKp7xJ0of9JpoxLmbIJWbDS5z0DYMyX
6A2L2WSazvkaSzAcmRX3ATtV1uXw4sqaxLBUq9vv/nzH/Rwo9u2rS+16ADQE1nrik/HxSZ6x3pE7
LsybVKCFmnnzTh7kuZuHFETSV1Fa1A7yuOhrwAOCWVrEZSz/M8DRU3/J9TQzfjq+HLneF7kV9zUR
7B9H6B0sEyhe/UxCM684KZhTPdWzlgGKS33U0l+Rtf+MGe8RLUO3We89/WCizAKMBvir5kQuQKKb
rLCTFYLSc1amKLPAbQ/vjCBXfzob//mZsAVELf8pseUHmpjhpH+gvg8ml8TdzoYBuvYQAqNHvIPJ
zg6rg/EuSmetwMMI4s83yFVf9OIGyERE5IAzdPk3kFbcYFMnbsrLMIWRRDy6IsKSLMNfZJlxDTsb
jSIQpM9QgR8tmRoPaYWSRJD/RXrL59Xtt/DsMfZGdDUDA7xxHNoEWpVYlQchjsgWi9k0WozvO+HB
9ZD/ny11jqG+tKk5dXlW5k8xwJ3oQzpap1SIq2kmjTSH44q6ypi6r6xRNX8Hccm0fNFC9+jbRkmA
ZBy0Vt6gdx1znRtVazuCb1Y5VsH98oYS+MdOwNB6IpJM2HJ5/eeTIZ1l8MXTDic0wHelVn9K3R4x
SjW6Xzs17RvwxvGSI1zsGEEvzuSS+fQwuKbwo+7dSuKOOFm+lQTsDG3DbOOvsDNux+4jhuzum6S/
yHYn/3Xs9ujl6xgUhVIAbdID9Iqz0WMTWpJgFj1zeiXqo5a4hTcnpRfWYRmxe3aUEbwn1z97Fr44
1gxP88/f0hUHZmUEDhBLC6CQCDhhtPxgMXaManpg4RdB8xZ2EN44V5yeVm+y1x5Ii+lMGx6bMD/F
OQUlGxnxd/FF4fjd0KRrcNjEXmEMCaFNcm//3/iFz35yFh5DGpHXa2RGHFRFS7KhHMmZS1CTm18K
KsEchppWzFArNpskO8U9mSnA96gOgdItr8LR5kk+thiheoxW2aKfdRsMaICRYZfnt/gnUdeukP5M
FGV3SEOMsZot0ZhuE3TBCRpYrk9hQhtWdQFy6VMLtOtRPShGYV9CNRxflS3XxG7TgukHvG59NyvP
P/8sOjNO3GBkaYHV9ondF+jog1Uhkez6t5ENIuXtsWwAZYpHHPiZC8WzQuzEYnCJIB6VHeYK9XKR
j0Zc02qQN9fLsarb42KekjEqe85asDXOPkZFi2C4ei/oV2nOTBb7y+4DCAzhGOoYon9g4lfX5cMU
cJ+yJzxqGvbS/sWHcAD4I5KmvwEhC0zPgTO9tORAloUUfTn9b2fC2hglRJ3t1EjlZSN9M63MKppt
lJk+Vv5T3mHpmATPIb49HHc9IJRIS0SGIiOZaC7qwMH9GzbPdhBrApoAi/X3FxKjr+8ClWaeV/o6
guTHqh3ATscFjW0WKt5JLHxVrvCG92bYwB74NEmmlm5Y+66SBM8OWBF+BtY2N3B0t5HSXtT9D9Mu
QAuQKxHDibk/7QLSbge95emg53uJe3dZu1HYSFf3kQR4LLiS5yppFshd6bHbqsp8juXHxh37CGiR
ZCTzeWxoeRLAeDcMj/eT3lean69o1GqUdbk6nkwyyBbfWdpL2EZaJhMILl2a+d/85iF8YR9Wa7og
E/MMWyWs6r59i2iT3SXwn4jz91zDQwKmDuD4zFC7AxQhcnjTqM50YyVHnxA4flKxlDGgNZwAjrL9
eeJGeTL14eQGJg3AiGCHbFngUohUXjXFKS1v8Ud1jY7ZL2mUbtn0+etSzc5kOfoH77m4Q5lJHnlD
bgiHrVa3AE64h43+WaNLjSnzGvUKoNO1vLBCQBpIOeBqHINtpuaQveef8SB/otPXmPwh0ZPQqILZ
QuUovjvedp/e76xr7C4b0f0u5m1Gtyh2cIGyhfD/zFDYPk8scx2cMreej7Npe4AEXUh+rwKphXO3
uJG46G7k0/VbJVQXvvtDTfi4H2qmFUAtlhHTiStuvPoc6wIoGkMRQ0nawOfiIPUaBqiQ1t+knfHQ
Q3lUV6jceZc9BLd2Q9WrBzgodxiv4kpgOzE1y+GjnbJ/Lozr3JY69o+2pGYVxFiA7+g5PpGynCHP
Uojt1Nyfu/B88N0ggdRw/DcUMcWkfe0Gnd1Tp1ebgx3UbDggwovBI7b3k5d10M7Zo+sM/i2lAGVA
0qujmgnksNBbx4YoCvJ9HdWvQaPMZtltQlK6DXRVg9egOKN2fn45LCIKeImOMNMo2xO9tjrnVcYb
hErPY/Sz1TvbTH4pVAhJNwkraYHru/SkCefw/oMB+gwMgFHKz/elGqPslYer24NFfGw9mg5hufph
oovgiuhExNRRnphLtn1O2yUcF3OmcIP4uHaUyxHAW+Cif5jOujZoy5vY6brpYHoPoLbcE3HGtq72
f9+m7s1IExrjQndqWx8mpKmsEcm4t1ss8naNk6Fe2tX5w4dai8tv/4eqh1yPin78Dv8r1jAs0f64
oZdoXKg9ZC+m/lAG3dTuToq/CvmNIxfKJ53HCeTulnd5IvT8ZMYhiDNz/HqHGwqIJ6R3JGm2g8i+
B/8yIu7zwiS9c7kLKScpXoEONXCrwUBBRc/7/U20sN1CqVbhRvtATeJ2vzcQML5DXRw1O7Bc2Npx
X88dr/KuIgY6Ba1q4HVsc7xTETMnRfSd9Qan7yMvcnG/iNx2596MKhFgEvSt5lJSf2mjLUux5ZHV
Czr3pkeQLQTq0Lb6/nO0H0L7PK1q4gA7AXrHa+gmfRlyLmskVldpT3GZOTg8+jQ71FjseY/YAAJK
CdsNo2rLggf5kcczubNgeZCl+TrEy5ZXb/I0Hpu2XXcfVv9JJiqZY88LnkqAtrRKxugcq44vqffm
9POnz5IpY3alUe2yDX+BVHpqwk1rGJw06FNq3clkJU6OrDrf0xqD7TR3H1fxN7mlODglFNrt35H9
GS4bckFSVcPdSVOky7q7BQU5gE6y8iXG8+a5/6dnqWe8yMaQ2kEpoKp9wU5gtUHbMVLoQYiICztF
ptc+ODKmybTR3m5HFi8bs/r+sa1hjNdzKCrQ8qQVNCK41pSxOIHf12Wt8lUkQjE6XNPT+dyTBHfG
EvWNZg/RAA05kak/D2Dskfc+UMQsuy+YWyw6yyEgi0oOss70fKYUIFc26dOI4iJc8/MQCczVlJPn
XCZdUDQnu8zMYZehQ3a1pxqlbN+ofiLf6ZUCG2tXa0eNOu8YRmDBJ6ykOc0n5Xg18rWq4Lxk6oa5
dv/05rBOGaxYUKcf3M8vuGVagq5SqtfG0lsuWiS4BNKp+sEKTuU9qU0m6XlMdYXBylQCirZKkn4k
0GokxQLkPReOfZ1PyxCFOILGBqfrVl4C769tuF8l9FH3UIE6mMGeRSYlujI0T/z4cXb21h2EePyn
MINDky2V0mHo4B6HXJqFoi2/34cHuDS740aO1lr0uiGpzb7RdAUi0S/yKwf2DxqeIvHTbAt3uprV
LdBq45LbCF0rSimc4ZNOQTnbNKTnufJ9ljbhHCX8azOKggAIMjRCj0s8Kmc1ZqiOiuvrlouwHHen
1lPYekshp/LjLp3i9o6T/AvBJUQtfxcgFYWtvKLLFFi9xLQysyFibMrKHMYvMEa0fWuy61KVH6y3
txTlBwj4i6F0Y/hofW3t4QfQSYn6M7yPZkWK7loBW3m3hbZahtJX6F5Kt05mlVtvFfKOeyTmNWsp
urgDRB98CVen446+KxDUsQy8I2xAisycHrJ2BHwrf8QCVQQ9o2n1Fepb/cifcU9k8DOGgJ0PwRcZ
CQP5WqAVjS2dhT2OimO4BP9pyoaX4YtsSIMFqIOvXr2Q+Ptbz595DGgtCw3h/wv2+NqIDXpP9y4C
LeowVf2B/tCB6Eh08ja82qFPpMzJq+reTz3rh61FufS1f4En0BoeCg8+LanhF3cjivxxrXOvO8dJ
DRALqCd+DtE8zWFyL999i0ZG2tzTyf69+M94AMFFF4m5aXYI/sRlK2Ts8vLUVdx5yCk+srwzQDJJ
K7slVBQ85ZeOl1tY9EeNxdlIMDY3Z9HOc43cz+H/zLdQW0e82k+lpiwQ/BkG2/fvB7axEaxJL6/p
PWYDIGUENjk8cHYQ9zI5J3BnOBU2OuXFzWMga8z92+uzTxx12NSqExL00iLwecXZnYI7/MPMaB2O
B11iJTY32TuPervqdjkPqSV09zL3tC/j9IwFpj+UUZ3sJeeQszb3g+C6quqqJblwwNKm9u0xt1a4
nuU9/OKeQwtKce2/De03pNRUIXdm+cXSQbrI6DYgTDaU2FNwxwVohHfBPrNeqH2mRmsTqzOSNAQ3
J+2OIpX04XI69j/cOPocl/XL6vOT311z9udOpCeODGLN0mj9y47MCAGgPIH4PMLf5jSOJ3pMOQjB
Rr03xTLNo69ebLuUZCOfm4WGCDSaMFsnWIB1p98EJjhuSRMgdMVlwTdOooR/0a6Sb6da1ydWcX0l
YOjXVOVZ2RjAnIZm9alOD9f5Fa8uVtDizhyzifxCbwOruhBn9J8B5jUmSva+e6oOIguLaLVZJCRV
+o3x+kBKgDNjrgYbXpfPerskauxGR+V3M7+IJdRXIAWmo1opfa/UhIjZyEGnAMwddXvVNYPcDp/N
22RXBjMVK8ASvJjPSpB7TS+blW/QplFnjXEaRGNc+i+OxQH4fFEYq70n+Ylnk04vY5tFW60FRy18
pgpT2zraXaC27nBwthfwIbKU54gEfiSLUmhWZFFsjwE15k/ql0UEExPt4iqvaPSvtkId1MFBba7S
XTHxMLhJsb0CJiTKOsHRtWfGI1agi4xl9jK3AXwmxTXluQBEuIGwQWAn9/92Ha4zQoeUtyAKDhWa
enZ9D/0FLAZ+k3wHNoNR6OsakvLjmppYPaCGbAZsH06aeKTBMmdNdVF35OI1nMl4pJ5LVEMWA5iI
ADPrYdX3xCL6bjBi6HBnKfZCRNT22z1xGAhCe/FT9zSppp7oFgJIouo3acFuNRzmRqucB5R7Kj0O
6r3VDoTBY1QHjndoesrxRAULs7lEYZSJllb2DhuI8u9LOYQFAoYgSq/a2Ss2T8P/EHfDrLJy+hSU
txL2K75ANljT8GIJp2ryuIjU3CqFmxLJs0wSJ1cJhqBX/E8JUE3EiQkqGimqkNlhCugDYOftSvhr
NvBMb4YYYiY7G62U+bZJZ6UDtOqFl4+oiVUtrLYOA7RM06dcd6Kxqjtktk8hQ5a/TZt5nI81qDSz
XvgKiSX5qE2+cDgoYntJOBAIE/OTsyYs4nyMD9OZYpyhd2edb1s7ILBl98Uy423P3b//X3MhGRYy
oDPhmIuQS2DSQm8yNRCpBbOpVHOb3ryETxCmxVvxf0Hf5lCYSB3Z9pqEuHP7Om1Ir/9AiwN86nP3
vm7GkTs7RrBxVQdQhVmMlSM84Z/oklW5DtoXJKddVnNhDpM0++tQo2bKPFpLguqkuG3PWWWVPoyC
Pzda5GP4aDADdI+KJHA7wHVgerqvoOSlSaJkSlt/Lqaa+9quSxqZoXK/h4d5Ly16W+vAeeq+XJKx
+fdsG44Rq0pwr8TgtaJ/Sdekl+Xg57dMsslqwbOg30DqfK8hBBSUR116KSCDQOGJELetBOB7n2cc
tTKjTysX77UA3CaROtOAuv/k/xK/1091EvRiuauTGzVIN1fcHiPWSBYBkOg3j5Y0uOGfkKiKhpUy
ZH7MjDBi8rVbmsVj4uK9JMwcqGeiuRyG7GM9L6+eLaKb8EI5RSuRNEv8CZjK68AoLUSLqtmvPEPG
UwmKGrFJt3eMLHbEelPZkTmRZ+4bFwF7pNL/mGC1d5v0xeg50lROkPemmCTiwtI2Qb2bfL6B5um9
vnCJuS4sC6smQxNf96Af+2nkkWq5PCHj45LfQMGWqmPgo3uBYeFVuL6ObtyV96qWUVGDG5ruJk9e
EFs6V48UobvQJrI82vuRTL4quo+jJscJd13aec2XIestuTsfA/y6R/DxQTI3sc2gu6KBuEa8dTx7
BVfQkXft/w4URcJhGlBEwzo+CbJ7VIJ7W4Ta0VRGh/AM4xdAE0N8bw8S4YaR3+cG8Ey07Vcia/xZ
VtOBT3u7E+O0uRkAg0d1Uud931XUHREMoN88Wxg/DqWGe9tFH5R2dnGQ6PJKvFtY8mXccCahtm6A
PUXzojEsaCc76kp5L6BQZeXAUiP1Uif8cB59xRqbb+KJONNbt1eVKuGNZ4ItbMNAWeCjMZbxbS3C
xjFzvVmaXDHhScD1sO6sTOoFB6oPqnaqcgOPgIhviY1RnWTp7leXx21oixPrLo+uEdSl38cAmLsU
L/KZI6kTAX++XMIwzOQzxXu2hpQVTkSBEsv5IcBlHfz+yHei2lDbqZE7h24pRVUHC59meBEtxw0R
d3UcWin/Sk8igdgNFr7QromBh9vOf1u0criQUon0b3kxel0KSVmJwDuyb/wNjPGtlfpVKhUPp6IT
t+5oMJJSolGvonRO58Kxm+ijXH9xQGWCrsLOG96EPMzbp0O+9v4WP1ROlKrbNUSa/WjzL390edpl
anNqcGk5XBpan4sXd5VETKxEtHMhxpJeq7qOqHy4gnXRCw0QBYRHZ/E+i8xOXrUDmnV2qFrvib/b
VjeWbTOt41uyyS6rbGgIJV6I0HR5dq8e0iW1Y82b67EqYk5LsKw4LjHVxf65qYsG7KWv6nJ8rzU9
oqNojv+XES1ehSntulqHyV/3vkwn0nE60z4HbRpDWB7qrlfHLpp2SwM47sJiufQgX1SduZLusfgn
4xHf3ytuaSGFHBXNrB9hH/oCPrtft+XPxJqSlGyvzTmorx6ZE08gDQylS1hkgCJp+HHp+pTXpQYj
RJh+lecvtqFI33nlXu8525sUKxT6LlHKsKQubczxFkmKmkcu/BK2L0hMmKncZHkEs3UQFBOuDpmG
uE6mHRmeAhTv59NbVMKehzCDiLlu/30DjkIP94jEUOAuW0o0oGSvze/esiECsl9CHlPzenY0tJ4e
qzMjyrUXS8rBiuJkV219jHaaiIbiBOEWcqvbhYv4lHioXkTDlxifEjiGmtrtNU/mfV7SZrA6d7Yt
ZdiCSV6gIaERc6ZfE3oMhwiXPtUM0san005LVdN7AgQLhrKsdjjJaMGJ7dtempzTGIq+3Uw5SF/o
0nyKHnuLxn00Y1UM/NZ9cwXi03Joacn1B6b2dX6oUFdU185IO+yDutAQsJae2aJv4hhBw76L1IGk
bK/jEW+kctL9bf8cD/tsiEuaNYeV5yHfvmqKSrXwEumlqUFLeKToSA3YqmSsqGyNW7dnFqlu4wzy
Ug7JIODXRE6d0m+YsmmVnFugLbv5+7fZvFMLWjcxl1aWh4+3MX+3bxEsVHE6D7n5XztbHE4e8te1
gCQ0IwWuNLJPYAsZwgYvQ+5QiyKWJGmxjcb26W643K6aI7dRkRh95shh0mnrzPOG+sSGZ5GJ5Zyi
LRrh27iotSAxBgB66zF8iUzaXGDpiFGmJhLGZnK9tw6aQ8PBT31J0GdiKP0UXovzQXbHcW7/xkpm
dhagW3rdRgBlzE72GM00N76JPW9pjQOJE+///OjxeM5oK8p4hHdKPXlDvek7e3o56ohmVxNw2JUW
q/IXtgbsshHkNgbUb1Wpg4BsdZ0R2AWCgk3qd7WFZ7ZTJ2uHOH2pXzLOtCjWI4I54OMdTmdl3YKH
T51tpP3Efiv/zmpIIwqaNa/2v3L/uNIML5KVMx9zrjwhydzkY3HSWyBwNGLjdZEYyNOm/0AZUbkL
tzOYWCeXTy2dWmC9erOEpzGTTlll1QR6H8VAQtRR5m/lh+jiXPK4S4ynpp3DdUiI+ylPcKZo5Ex+
q/9sE4pNS7MHQOnQYEMbXg5leNzsxRNEi0n4LeGY34AMdSwQ9Of4HpgrrX2j5bR7Cicp+N1584Cf
zmWpSlE/JyYhYMoYOVAZsiMhxvSInwUHyImDeqGO9PRHjSJm9wtb03AwDfJ8oIiSkUtu2xLIasHf
5l/9JxyHknQPM+MVEAmkD4iFX9h3+Dknhl8bGQjFLMloBUYy119GXd0J/dd+U8YW42OKrZivSUBc
37adagwoy3G+/lwssVTnd6IbH78dwrCTLTVNm/DsfSyfawMYt4j/vVJDhk9+H32DfXQErBBHEpEF
9NIL7Emrkr3MNs8sDDGXlbkQ3vSAR1aAB0mfPfiLBgXPU3cg0nsIqkJwsrqVmvm44imRqO9Vutl4
KGQ8NhuMDmaGRfwMz+9a/xuARP3BNx/nqeNbY4R86ugZ6SLl+jLId0eRg5m8jhogxasps7DGOyVa
zts1nDLgELhM1EkTQZsuscM1mgiBDZlZ/L3Snqnnrdufnm/AVl7GkAmEC98lWzdNCLT2Ibdb2YED
NV/vEStvWpQoZ4G5XzeGvZUUsdidSgiH4JcPxQ8IHAEuNds6AvdOKu5JHnQA9kiW0kXXVdQWEy1Q
75Z74Y9JXEWfBKF1PdWxjZdUGdPSaLjbsSKytuQUYU9CYvGu1VlrU1DpsEJSFgDYr4Ii+8nR7anD
/Rnzd0Ovb0iTiMMa3yVqpANAozbw+sJp3/7JjCOXEuL1g/huoydWV6bAZIqEO9u7kn4zsKiqtiwj
1XThWVseC1D32MPAOCaM+uup0jcAmtc+p7BHQVos5WJBrK1GXCRa8qMSEhMcXS4ZrheQVyT0np0y
PEOZviFqES4i0HZW1EgJ2rDA1plKeS2ZOQIQOeV29daEx1YRuz4Lhfju0ThFSNN4VvVb4TrblaqN
dadxxh7MKMksCL+huAmAfZwhjw1kICakG/8TXHWEgmamUWksaeV4/X3lIHZERHKN0JVZx6CPzTOs
+lu6wimnIaDvWnTnMw4U/cYtJmz+eV1MmZepJZb5ue5IahLSAijLRb5qg0bFGp04W1Ksa/DOwmbg
fK1Ppj+pHSgv6OtomqHuh2cZ7QepUC7EVTKqBxvyQdgOxlVf+LdYYBm2HUML6k/jEtC415CXmR0h
RqnERfj4uDQ2c9aILmasKKxKWTget0sA6zaOlG6d65oO28hXD9Giu800lECx8Gwp95XEFrXv0EZL
Z9+vZex5KpASj8as3mBHPnGFmrbDQ0JKpbHWEOcMxqifWqiQOAZNPb6aSjmO5mkPfmRJQ2W3GWo2
bgLeoerET/5BFBIq7cf1gwo7KtqDna66PK1LD6MJqewtBQNfhjOVePUno4bRe99Hj8v2X8sFQdox
mXZVIxZot9CrlUkRB5GAKY8thro42XQ706vgqG6K6iCltPFdQlpyeSpaEaBIvJPFJPyy1T4X0IqB
nREjfE6LgJi0seZQ/0FtHDl9NFqTDjTW1u7xztzK2LXVrYvZsJ/U+9tYUZQw4Gz4XNknm4rq/MKo
YBq+MRSa7V+KZ0mNneYvom1w3u5qLep5kZuNH2cK4eFEgX9chSErkUFWjzBVnpGnr6SpZtap7Hs4
Sl8+f3u2drHFaLlg4f+7qZAArY4CQ2D/X4b+t3870gC/eEM3Valsrisy+c8PaSkgmJuV9cHJc44F
xrpQ5x3LWTQR7EqVnOM7ffrOZUEVVT+iL4LPn/joJ8WQZknHCjSCDBNvGBLnNfVju6hRaYimUX2a
0ViQ1Kcg4c32QVJeiss9aeKTzqy+VQuSdp7Fn7CFcbKAhEd7Ew7xilZVRSkm3e92syTHYSFF02sK
pd58TaV2+LKDVpDW5j3ip58waKIH4GtkgZYkjKTSaRF1WpsnSRKSFczccbLaEAO/5MbKAAUsFScx
WaeaWJQFUL8BjEM8nOu2j3vFshlHq/g42qeeg9axqCvnMLr/anW/CP9Ib8WaG3Jo4e4Rd9wq8Rru
KPSx3vTF+hJ6s+SEZFXS6YWBQ+WMv8goQ8cF8mkl4DY0uewt5wtYFam1e16ieo1OjOrl0IEobis0
brioxx9nhNW3DzoBbLGwlugApvcnMQegDFo4lR7HFM0y9UZ0rRcxjOemPvB7K+AEt2tZhPCGWURH
UzAavJXCafpOZzwhDYI/rUm7p4lQq+fitEsAcUIy06C4BmLHEJB2+7cS/QPZffLz8rD+tQ0z1c/4
e0dBAoZ8BeqdUMRzrGpXTwPcFOI4YdcoykNhBcPjbqlGREH4jDoKfkj4fPqphaQMi+p8H3PrPcG4
wSBn6Febxt1ZVI+E/8g+5RWh2DxtshoS8t/vrkejPA13tOgYf/qXS2Oyb+77UH4hwt5XGB1FPRTJ
gKpXpjbX2K+URlhlCX66l9XPg80sGyNsXHbctwIBiUmm39wEukMbofwxTNA8v75/vAsVN3laFAls
rr2re82CQO+yBVXPSp2wMACyPgUXDpSwodK5+Qul1B9UKDDPsFUDxeDqsdjenW3NSYEZeqnTFNgU
A8SM4yb8ru68Y+6ovOIQ7s5EYlXw6yVOo1mXrKRRiT89oceuLqohHZWmzk2c3UwBaly5C89MLTa3
Uhv1GPwI0syHEsQrcK4cgeJBtKlsZ0uHGyGBLXlexxni20HjWmeC0Ln2PMNLnCGDDAilrAedaBiA
oTm60XBCoIGaG9Br3OAwBtNkTEL+nHSNC9kJlANAWrcMyc3GKUrYMebBI9BoG4Lvn3+jnnM5ox8W
e+nf3YksqekQBwvIrUsj2o+XSMBHwJ3zlXg/PkjNkGDDm1lOPd8RYpas5HSRIOikymJYkJzJBIJr
8uz7qJeuadqcWfGQhZkupiJ8Oo/uYbjPM1nhtIEx/xJGK1BUKw8w2IET/5Vy6ZSsdlk0JNvM0g5P
nzFnd3TUwkccUIu38Ek5FaHoNqdm5TJcPkp7NeCLcw4Jv2URXj87delm+UDTGrebYU0Ni3hI90T0
YmUDKpXjcUH/lJJay+dfJ++ucZKCvvX6op52tlCrTaf9cEimjELiwQwS4nJ4gWGcbcZPOIT05KKv
UC6YYdlfFljGBrU78xmS6yYQTj/Uw03qnXmnf7xdEjddAkqIUmxgSxb+yzLprVLTPi2W9S5Yegdn
PmiRFWEUR5GpUNIzLL6fqWQrvhB+n7W78QvJnAYGr05eUrrwcXKk2SetJ+JkNMkHJ1KE5c368R+l
NvSxWcGAJw8hr3dsJnv1xuBSotHK4QUJugSUqnHT3R9M7yR390GN67A4BNWk4JEzDRYPdw5hQSfC
rj0VEjp7zG/w7y8PY9d9VmzxXH9/EyXemV7QRNQPRcyHyKchR0nTx8T6IEjJ+YOpifu8n4PdPqXl
Gy2ct6UEn2OEQAWkhHsudsUXFVI5SO3k7SR95jeGMEisE9p5cGWW0fxRU1/+UFuliZ5xtYHYnZIU
P8UySdkwKp82WhpHtas/br/NANGh82EfON2eGcUbwkddk+unpS9phShkZEPxJuLshSkPkB4ciOGq
bKHEKCned8n3HjSUciD0/ZRXPiXDWwK9f30owAUY2zNpXA/7ahTkGHsjb82P0jjQpH3Zk73T99j4
5EpHOlSPzaeSS9X1XaVdqs7xIogzp44/BF7dHztxBwN0wQx8iEhHJc87rR3Y9BhvkpwEEZ7fnw2w
PVqQ4SfjFCjXH3GDWh3QEs7UTndUKEDI9O+xOVMx0D68sNGF0RHpV5fYdG3CHe3AVgHwbi0ofa0N
XjxoadgMp0kRwlyp+lZ3LDsqgD6+J/aA5Fxg3n0NYYxb8ALCfnu+vCsUxWPWFbMAVOT+5Ym63ALo
Ge9wAJAN3woc3fpPRtK4uSSQ/V2GoHbuinmpmyw3/3mzBOSc5wbEfNY/Raqbw/pQ8qmBubE6vSLx
KBO9/oDnsHaqwAzA83A0ImO54r+ftEnlkUsPLwuxwRiKLUCH0eNOH/Qy+zK2Xci3AeuRIC9qCPx6
wFZqT3XiWdSLd2BpR2the39UMq3GsU5ycOd3vHcskQXKh4YLYMBp1pyM8pX2Y3Yi1ETCMeH0mPA5
TjUCWd00ur5mxbCEkQNKcfZyZp1UZ0BwuBs9f85m580zBEMy1xK3zewX/9ECTHbWVzpFG4N/ZQL/
YGj6UNezLPddRaWA9ZBsNZDPaX1ZqVXct7+8YZgz9dz7eJjCmCUqFcL7aA5bp8ylDNqn+rb8JMHa
YpkKubyUOxYybY7DEZCpWDN9dIby34HlnMK6d/qs3QI+6qdoweKQD63IxSzVQdRBnBE7HbNTmjQN
a/5Cmbrs9yDbSzHDVexm0OVAQaSjAcEZru692nqWv+aisj9uVV/SkFZhZVSt7NrgW+GoYxJvGu3i
hVUMj7qcaeNWHuuQr6T5NVZ0BQ5iEMmgcLcRclwnKBdqJNeLkom0Yw6JgE2AdGjMkR2xmZfgGPZp
C2AdqvkqXnFO7Kz34PXJOWdTqHbXC8x+wvd+N+7QXpMgk5//lKtd9ckdFYL4NECc4wsHH0IHmKn7
TfsYE7EeIH5GOpCjJezZYISH1UiKWv9qEzF2+4zoe3xzIvQvANt/aGiAFAUUp8/jyW0MWFUYJJCt
ZX21ZhKKWg1DFaGyixfxz2VFO15opQkvJX7O8Icihx9dKYq2JCBoPLTwQaa/bwhVjBPw7tjC/FU4
/WHt4DiVH2CS/9KBTABUNgSEerqVggpv+ZVjfT+UQo7dnK2tlTCh85HPAx6n5mYLp4QN81GjDyoa
8RciUpjfHPBPn1KVTZgOE2fKl5lLSuqIQNl1DaHNc36I68M07RRG8+WujmVuk6eame26PE3vsWYB
orXRPzfy+bJ6pD5iCDvpVs6OcyMX1rL1VTRNi/cPRz6KkRJfwZCXcDFqJLbGwhnukq++s9XEQBBY
SrhwoKJHrI8qoXAE0xhgQH2HptY+X2awmtp0TNhet+yvCYe67ALllGp3+gppwbwxqw61jb98jb3G
BQZYisgbkhFav/+Ud++f2Gdg0ynSzHRC5iQA8qMvvSNtc007QOAsbrsEOqplnXlz3zBNoNDnfZ86
LUnwyZt2HvX3BlhkPsbXjMCr6tdGPVsMWaWNyHAbO9EoYWeJz7LVTe07GpK/ERQ/ZfxMP+kurRiz
pNrssYb3271+iVXEFQZRQ1uhJzqQOtQqeqdomZGicy1+GJ8OHLdG5kgBAw0mSCtz8uWdm9dwlTuB
/8zvjh5aqPBzkENwKNHxmhjfgSqozWJHchcR5Mu8UPQqsgQjeIGgY3QopDwb+qfxExAwgkRNuWeb
vm42sFLTzmlqh+YPKXGvyeNrykg2Q3EtPIBWe4qlfWvCmOPMsGmx+Se36BDtBYjz/PRusrlJRS9I
rSl2nssanU6WwtBdLzGU0a20KPo+W6LCmp2BQo0xJ5vbEk2VyWqoL12/VllZM1GG/2LCHXGXqIRd
lt1UVhf7U/txmBm2fJ40IVzKqzilZsTUM4w/Fw/keGIyzaPRR4I5PA21mcAgvqLoz2h+fb/Ne0te
fk9hQUCML07Vc2IhrKzqye96cK2QV8mCWr63wa8HX1yUDCLxU5bwzeX2yMnug+x+rGMmKOFmkyzF
+uGO6Q34bY2Qeasfu4dlXoiR2aw806X71WHpBAxYpss2NWbREXaTgGh0rog0jvIpOWxXcR1eUARw
DeiV2MFmKT751tAdhCB5gw/kxO+9qaSnVWwhA+DBXNbo0txDRaCG6dyPY10XUIrJmwKZ84mjMVyp
xHnmoEE5IMUOBq4qi74knQSF9MkKDmjVFMvhcoBUzoOOnPKzmJJohz9KFq4qwWucWZI6VUfnXcbi
n7gdATZLP3dXXn7gHFO4K9IcZDyZ7HqkMFPjbyoKj8rF4IAwIHrZlWVv5mY/IfUlIvunmda/Y3zO
ynqB5cUCP4XucJEyag3BvNa9vFVDKd7426MpOw9VXe4DXxyWfMaNIwNRCbnyq2JF6JkujTCe85I1
3htYxE1J3nFQSsgpaeeAoKy2PwdxthYiNMdelByUMxxHXL7wfgHLUcqCkCiF5suWYRO3uTqzrJOK
LztnOG9AeIFMLi6m9cNjRd4Sk9PmiAMItk7OlzFPi3nepkeYxMZfiHLzXIQiyyVWS3Y6wFM2UsrS
PmJS1snF4dojq/mi5XINDLwm21rpGh9KwkQR6H0/9aYmKZ1PgYM1o9W4g9d7guiLFw2IvZXeHhsO
KPoMozTaRzpoe1uMWn5dTWlZiV1rbqg2ZGIH9EGi7k5iMrbU7CTJxu4rwZJ3+q+GZUZQVihsGtyV
nJPEO6iwsJUgPFhThyMxh/LjLYwDPqrQ5bvqLYiJrFMSbzFwkZzoMSvkuovoBzc4Ymo7CfhjAJ4w
p/ljRfSOeX/Vv68PjqHllL0gAcy6hB8bShMO5f3ZQkJdSVwMNyBEQSw9GF8Wi7r4ji/64pltuCzH
mCWl5suM+cEgr2P/Vlx8oqgUuWY8zoAXj9rFnnp8K7Cd3o00OqbCsqPBjeq55wAE2HHH/ECULBoh
fsNXCDVshq3XMoUS75tfr6I/MLwseKePpZL8gG/DzZaIlPJ901P0c7L62hPRoLXLkH9Rxsfqc9zy
CI2qoqk+k2iWDxlAM1Ci7KAlwqfHs4s4v9MrEgUHlJ7zirJtO7m18MgKdZIAVbYCjggkV/6d9KjG
PeCDI7hm9KNM5buz4qdslQcuV6pHdlIuT/h7tDFND2YU0G4mIxkzg2e+zHu2I9l7yoWjhrw7Oet7
yUALAr7ghk9rZAJqMqpzvBSO6Fb58OMK2hOv3mQb9Q2hz7F4BekHFsusg5xcGor7P9qpwtobGMUk
Tck7pkec+VeLvRoDXQ7BfkW/tz43YRc2mV1Ocr8Ekud7Kwt48qrjAZtblNEblFQplcVbPB5ZwfN3
SW6gu0nqr23XTz1DuKXVkK8dZuSTNN59noQqkWBOKGWOk2msH3IQSush7AUIQxfvuZs5BdNL7J80
OViGVkLjVKihZER+jiEJlvlwrz4SIdYVzYwGcjlcjKJWXGQH4RL34H7RF9dhdzmfyyxKMdW0kaPs
hT8K7mS5u3fcYN6gnXKPa8T2u6eQWPSXl8xse6A3EC6J092dqZgGqsGbpDtRg5fbdgNtXl65Sra/
gzDsQbzg89sEuakFG8Lvb0o5D9pqg3Pc6tp8cPG0ahNZihO09bd4j/KYCM9nHXy5ZeiPHtSkU/Ek
bNc1/n6EsBPWuQRLuWKgkHDS4do+nelKZvKUrWCd9QupYUwn7YkJ7pU8CPsn4YC5w57GcGs+aW0t
Xlbijgx148lDSn3BUSKKLE9prC+Ww23UWwBJ9TJp3Eu9Zt/p1wMl5jxDn9ChI4GkYqKNWm01FclX
fUat5tofSNRu6DHoaKGpLKt9xJ33GjSwigsX/7b71DH/6AwIu0Q2YZgg24sSEY/hWn4DwXhX5SHH
MUCXBj4+fqbZwt25Z6KSZp85dHQxS1RSIc7+M69TmlN1X3T3dw1Z2yC1CuHCy4wZvoM7F/NxBgbL
1OQhBiSCQ2NRpTJ+I4tzv07NrXaIZvWcmKZJHxmlmW76uYkNTAYycda77mP3r72xH+4b7bMsG2ND
eHf7l1YodLUU8131v7bAHWdND6CbzeaO/knVtl1UjrgiMWsMWW+uGku7LWNEJFLS6Aj5EEZvD9mZ
aM/3bBzhFGd5STBESLdd1/VXyebKBAlZc0uZSD/9Vy79JOfedRoNe8fhMWgNlASGkNdn2KoKAWSl
/zP4zJXIOXCZu7O1TJTtM8D2B7UEdfOudV/HvCYjd/SiDl5aChiT5m7rq1hgqSKmtR0B4AHIwXMq
b1ZMJvl9ofhIHRH0sqXNU1ea+mikmaadQQ1r+Fm5jVqZ8zLm6OA/qHm9H6R470m6iWGkminBmiSY
9IihpzIuqbrmVaCmiS5sWynjns4aXGpDpOAVO/bi/XtQ38IkxTbmj5864WE1zP6R4VbmqgLDSOaO
GJUC9xhMZNydDPFPGEEEBtClC/sPcQQ+rOIPkYc//4v2gegUX7WqUuhNgZtRgbsq+901VJ9wi0N/
N/q26Y9bamTGoQkyK0geGCi2Q037Lp+M6jnPZBTSkCJTa5J/U5abSgfKkN5NxUjDNhMkfXxWc32x
H8I/fv6VBRPrenInjFmPyyijCuolbecgs5+/9/R9pcwYC2IAVbHLMwCpojx+mivNwxDT7IObKQD2
PVvEK3eCSZZROY1VdFv/bqf99ZT+q3A1LXkDtnrWjS1sulokNJFG2d7WFstxoDa2+USPvINvf4Oy
3jl01rYkr0Rb+FFaPNtSnSoC0p+IGZrXAyeTdtu3oVICwBqVFTpfu/bZ1QQV5o7JL0UCrsWUer6D
fLAPOzE/OuQ/FokplOQlo09v/kb8bVsLhi2JRWWh7DCwLaALySekSfHlo1UK45xPOTR6Sz6Q1q1D
UhWAmCXyWh8AuBRTE9sj7u8ZQKj3X3b8HyA0JhL3jgqM1rwH2XTcoyLZgUS3/u53TZxjFLFvLGWL
NaL+qrSpQb8qksKYoMm9uNWg7hmE0H0SjD/IlQtEOwA0yzH3YXl7PLS3w+9WBJc9oYR3gLLCjvZN
A1vCSZMzTP6cVm7/TOTfWDiNWiNM+ZDN/WdQJZGGPjxzO+BmiEhHu+2FIr50aSTyeeKJ5LkY5u8D
hTHLSK1JCPi6MJQe4FJwR9bMnbByYgrDTF4Et0zJbvdlwRYRIOOntAHPw4Ek/4GwGAYnfmhJK5v+
yX4K2G8dSCFUvF0OV4phgtcMUpbEMWlMGmXpQTuAwI45KZTHdv99Ag1a6YhaXlumJ1L4cJI+qwkD
IHeQX69Hj4esFqQvu17mJ6v8dG7atfd7DwxqiNHtiwVkYyNdPNH8ieO08xxa0vlDwvzdbWu8sDA3
bU/glPSoMHLSHrmrXXPDj8pz6r8RyYrycBYPMcL64dkdV9y1FOTcDgng/HAI5RtDerLqluYvw5V4
6JO63JqmvR1kKDRYp5BYay7XVT7QktaALoPl3luP6eee2zKBlUHctlT8hf/08Mbwt4b45EX1nxu2
a4Y1Q87KPT3wvf1q/Z5Ey8JMRonIOzv2wVX0d7W5kz8twF7KVXjvipRBvUiTNsPCwr+/HC8xMpND
vtzYPYx4LKvx+7zU5ZgbaPeUJ/CV7/Ltb5h7LhSgmrZa8eIhNvNoiziKzwMoaN8rNSwVPRMeXpHW
gjegatNOM1/VFq3gLbLyZcZQnl9zIVcEUf42o6ZadljfG8CBFGOsAfulbsr60aWKTeMctC+3fMET
30biJVVKDq9Y4G9pg8lNES7AcRUg3TkNNamf3+QlbZL0QZ83QzaNglChPqj8PiVjraMkmVKmC5sp
Wm7WsCuGV5FLCHvNkRSb5h03MvuBHGgf2fMGYlux+IVXxCSpf+lEm+lfxC9JKm+sCvhbH1IERnlh
agEGtqApRvuykqHFwBX5NyqFfxjzbhYn2daqKTkWS1FNOHnAM1GeteGYqs2M+ZDkUGPUGSxqZmNF
vR/WMFmYKwVHipkicPln3uf9guTG2zaKdpKS3TbxSJGbIndJe0LpJimc6aXkwagauAzzksCM3lW4
4nS/0A+VMlJJ71AYV0Y6wrSvhN/8DL6tOoOjWcAikfJP73Gynnvv4Q7k1MB1NgO7ei7l3zrOrTTG
8QIcjiPkyYT/Cpk1h8h57CqMBZXxK/Pk8T1IRjzZEPDydEwWwApyt8O9TH3k5dRiskxe1c2Ksj1s
L5vnfwJoeHNlZnFuGInOpPllXhSUgL0vvmlmHvvYh9rtMZ7eyWRknSNe5fZJ0sPGJLMZfEAc+DcG
iPx95vjZCERcxHI7m6psW2HzXmP9LQLApcu3OM2DgHOE1SBRyBuS5+BzEu+vV+y7VhLQT5UAf8ie
i9IeXnxBWBTZb+07+KWmWoUO2RnvTUPcbMiw4FzAvs6UPkZpzKz81XskwqUumjggYmPt/ulMCQco
/ROL5v3si9gSTYMgl3j58av24+iC6JeaFaeogbFQhRDkirexO7qVyCqkOEnVeAdGwstt/wZ+6lAk
OwfeFHLlnhUeg7hq1YzeXXjqxFgw3eT4MzHlAyoG6A56l0b65VJyNXiHKh2T/mbVFDBlkvYhTgXc
DUSvIkRwqsmP27CNz5VnAlFCLRwxDIJRb/fMmGGl1fyBYSSgio0UhSFUxYdNfdT3PXhZGrfTod8R
iZm1SNdn6vc5j4LVMoVqMbsQRhKd/jqtgpAHH8y7Rgb69rK5XCMTZgv1u8C6L3ApvAIWHGfLh+Qj
5fJT1klrta8PvtEZRAai+dxE0KblUG0BuEpz31MXXM5jP0igRzBYY5AqypRxOkBMN904UcXfSpPB
g+agesxw27WyCDCITYK76jTsQmPHVEEN0e7AOHcqtOPnbuFJ7cqZPPNcFqvLhVjfWyINHI0VaJ/a
9zQN8J9PU+CfAFijHDW/Utr4QPhZbzaxgNUdlyEp5geyC5IyOxzfJGm0cFASf7RrVPTLARMbAwR4
inpehe2zXK9/gBis79YJftWpGqo8zu2nuUaGecZqxQLNys4ZcZMdN0qzD+Bc6bqfft0TTCgHRNq+
BHOKx/Ba2Rh+WA/osqCTtUYY+jGUjRTFE3FLUIjMJuh1i3gCsLENathGj6tzcBpDNRbWtUyjs6g5
aIqGdxx9wIOpQdGvFN8lovIQimcyKZoOTL20HiqEHu06nMCACNAmwgXL8LG4raNnNRWGFVxbGYgH
Icwk8Khqd8p+hJmjOG/Ar96NmqffdglPthdnWHF4IszM+oTqPzd2RQ3Uu/pmCsYZ0LOrBPoUVH3J
do5NYsqujNXYO90ySr708X3suGAu3QqoxAj1kXiMXLrxyBHCK7+PJVRxWenGbV72uei8SnD2aXyc
xHpkC47FYYHR3OyMGzpnsRF9/SAM74jxUg7C78S1ePiu4iywzzzzkIEoinndwVb0BQoKuXxNI2/u
dKEuCKbKfYbWEqFTzk/IS749oWtb1mViQ9mOsgWl2m2LoEb0TnwpYtMovAkKg8VTdXabdVCmLsrA
ctR2FnXUUhz7laSU/FHXG1BqZVqxxRfqTuZjlF757XWBwh7rL3W8a2ODjRPcbHCfjcvmRyHvn17V
ODYjYTqfm+sbCCWTMoWzPSjpJaW6Ih6404ziEC/6r8cMEA9J8l7jPA3ZsIgvnbuXItwl91U0ctW7
yFj4LeVDAjMeuAqacmGZNHSKDM17QmKnEKdA63wjkUsT+JrhuoAYoS9QFJlemE85jJhNohDuvF4u
IiFcSWQ9NR6krfYxqlLRPc2gciLIPIbufHY3d7iP1WXzuJ6vJD3s6e3eM5xUS9i7qAjWLd9AodpT
8i1Ho6Wz4MXWqgbOhQOO5sASmmV8oFlCkglV6AKqPhimkno8iQ4OwASUpNdXYsztbP8gMEtaCJVX
RKkfW4ojFtKy0d/PDR3TbDTU2e0tCMbFg8yy3ggbGI7oyKbjrzB8DLZee3zz9c0jMEgkn3dWkVZd
RBjmeYHFEh4Zawoymj5bNhQeo/W4H4bCVzpwEdjHcqGolxP2WIGqRhdDLayXWIXGmXsb2Ho2lgbk
wjTrHdJ0gZ8BtgREV0q9eDEO8C6PzITWSyEG6WiDK/reLx3DP9E7HwLlf5pQO9T87qI3ucsk2Fux
eNXqMVHfll50JkSRmENWn9IhRCmafKLrNkV/BmmxDKq+tAHXPZNS4CmeZDDgufSqjyN9kCyj6xWw
W9dG0WCrU3/Oce+ahZ7asK0AzFU9raK7jyGj+Vtxw5BL0cx6HaisvO6rj6YReBlbYzCT/mmm9bgg
qvG1IFB59B96vmzMtUx/qbcYj0TQCvmSrjh/Vjgkz6rmbQfYy1oywOMEOAU0g4gXaHHQpSDZLhcq
PwWlWB1USfYUWLokrMMPTkM6T8QrvlkAaG8aVqrdB+SOLtzo+RSmqmDeHUK3ioiVgVA39zcxoQOt
kLMlRnGrfgCmTWIS0fu3prSK01QJX/RVAuEqGD2/oe5xpgCnBiRqTr9qvm8A4HC17RBkSTq3YjdF
iyQ2j9saP0rMlLfsWBhIsxD6cHYgb9wLIItUv0Ww+W3MvyP+XxL6V5I2QxL/ObrXc5zsl8kQBbnm
8T9MyB8OG3W/zZiO2BW9cDlgGpuQ62ntzdbyDP3oTbU2wI97Fw7QSZ1rFI4mS56YGo0kLGAlrr39
GvmNBwWJdlJwxt5BY/gTngvs46BpOsGFoJZnxGPxkWfsWIs9HsIsv98CpetyCTcd9WuYQlMwh2AT
JsMGGe/i8PNl4pFv8gdO+uxRc9Tm06PQr/v5wYQPnYAVlG1vgtQNvfAjV96VNmYK0hjNpTlLqz2y
/hJisQxIuWc+7czqXLUt8rczKWEuljwm/y8LgYUiNNZrr2Yt8MwoZ0pHrYg8cEYCpmuCoKSi/ULr
UtZq5reOnrnRibf4ISY6l0qmjDzFBCNW0SYvsHv+jfEG0wW6BVscTyFfz3qYTADLQ2vnpZwN1Pjp
LJyRjU4ryDglvTW6FiA96EmfRHCH35G3l0jI+VdGsA+Sy05bcjMuZUXXspLvxqDA8weUkeWsF4R3
hRinIzJY7CPs3KXZkvs/DhhKwG3FpZnKpIg4S4K8lJQF3kgsT4S+tn1nywZ/LMDHlXDC/tN46izG
Zr5xfDJP3HXwVoErNHEvyGEotlvn1/yPVWLcmmErtN6NdXevhNdMGiYJQ+k2Ir4j8l1DXcZIJfQ1
RJ45vl0UiQ0gkpIT/7wc6Cw8Lm981LiGw+1SJX6DcOB6hcLLMpuJWQpbF8lO3/9b3LrMoaJJKPiU
RMDVhOhyaV7Ly2wMIdyLywB24lCzE/b+aXzJP9CNtyOKLE2Nhb8nTgu56TEKyrVjALLLXK8gj8gS
mYFH2X9iUu8BVNFLDnsKaM98a+fshRb8rc20CCJzYDgRasLXqcR3tezwi+HgOyseMDtNlb9Y3Clt
s/yCDQq5K82yIrSzc7DmpZZatP/vbjcFZe2unPvU+062SFrvZeLz8TGX8dZkGUZySpZu9yC31phg
AgpqnimfQrez+Pz1UeG0MwKociC0H/4kOAdIAXx3eDbO2UYULFdzXDvDcLxE6+aft4sqNc/6rF3c
RouLByUZG2eDtCMzdUyhBMMkBShaK6EsMHEFvNZ97AGH8zgsrJkgBu1y4c1PphLAZ66BJmbeZHoE
55RXr3u5qmoA8D5pEIktrsEQAKF7Wwxa6xFF6VEdgT3izbej9tqTeKjJHOiTksFlgEBpHBrF55k1
reg5xBCOL4kKw2lQ+wcKycTmjXlebhjx03uljxHEEPczEGI2FtbXk1euO/LG9IF+OuSiQXjHp+jW
xqSRP0wtLE/pqu/mdgCVUeHziIBKt2eszxwdapc2tdqprnRp2FkYKAVB7YkQoYLsYu+/NmuetlML
GxjkV/TA8ln2QwdqiBXV3r1sIQ2yvt8oheOBrrD1unJXEidDKT0HPRF+uQjuJ4nGH0Uo+pivURqJ
GqvRTYrwzyu7aNs0RdZloS5PeCug/yOSQJjBW/Ht7WZrUP0bGqQzYQwc6VLEhpa0kRCJqQ2CMEAr
O1KhsebmGGUAP0D3rECNL+po7s3PHQWN4YWcTKUpWU0oDUJUUMPNBCNkwynARunIO7IOrCr/623P
3CFgul6J1wNflfzHOqDTRYTw3Xip9HakRbmFrupxS8a/nldPEU6xfmprAS74Fvsod+rlSXhORxzy
uD7ZvDjtifPxmLR8PeUQoCFq2z+wgYrqU+g5CvFB9VCdUBRsamuSMCfywtnH+BrseGLcuf2yXvaV
0tDqI0F97JyGJ6kurkmAMeBL6fnu8AXxr/Qe0xmRSyphGvWrzaQuZWnv07kGvd/ElRG0/yzlxjMZ
bk0jWnuu1OJRH4D3j57dj2hHJhGaHNqnp+XJK8xlqoabKKBtjX/h2meL6WuymM7u8koA/bNsLOGN
DhJ6TXmITexny5MQYyAvcNCLqSD0mu0i+Gcq8bTpGBpXx92cdGD6R87UircR6bkMuG/x5vWFwFrF
Y+r6AUqkSlUWjwBpqR3aw1w+dsv7fUmanFrzh+m32k3Yn9NM0GE3fM/LmDZFeGR3jodBFNyuBDrl
v0orYY1IuP4cf+d7UM+WVOVfUYPei7h8uV5mjOYobQw+u2+8p55my+34cKFHnEW37cpA4eXJOcOU
GXCpfGB77BbfWGNJv1+Y4qMCfDYtJcMAFeWo8GeLZuisGOyva88NLNAoHNT+rKYAVLnTqcqHM+TC
BWAlKxax9zNKDI7X7gqfTPTCYP43/LMgRTrnbVBf1nwZxAeHso0NwmzeIc/cGHX+A7eRHhbaER06
O9scAMbZkVqKa37STZHV1cUSaKXotGPncxtOPmC14naLw1RuI/5R8+f794X2wuV0RkTzSoYFCk1S
QV8Ngg4gmd4pxaGpxPgECJ2C9AgVmOJ+f1B9eZiTqLwi2m4uJqSpcxiYNX7J8ejzkkDIDjVqD2Mq
aHU5GgkwJr8Mc5f4L0mkspKUsxesxYILIRDP1dN3HvHx6crgwA6jPs08NhoUbrKrBkDYPODHNQ9n
tFZA6FQ3Jnf0XKxB3h1V4khCEZOJkFSbkG52CGMWrvqlnZHNI2pKy0AsyDWgoRtWQcjd5XLIy0a3
lN6nCmzzBhbbmg7PpB4iNM1C+cE+u4yCrMiLQdLPR5s6KWBjuan/hb6zS/+lVdnNA9c+Qbekd0i1
x92hwlB5jlHUfmw6zFkpEwLTUtmRTBjAp0+Ixkt10wT3wOG+N33skv7u1Vzq7/eOqYjsulmu0J8J
zFh98UrOOkkXCFwpH2rXJCuzCJKpcH35C6Uc1GO2yQuMqHwRzHf1xxXHHQwvb/mYOvAXNw9EToAw
An1LTROMua8Lyv9aMd+pG2oyrPadHzfhz7ndqGppA/L6wSZhoHfdcIC7o9nF8J4J2RGiWTBXGZYr
8yRRdp3oKA+/xZx9A18U9+KIUTUM7vBYeAtA+b4fkqW1x4+Pngq8S3UWlMcukHEdBj4yt9hftGHt
JqJIiwKwfix9RPYwvL2XN9+2nItXL1Zwbfs81+NCL4ytsJdbVNsJGsFYNuVncQ0tUT07Ns6QwlBO
XiRa7GKXW1DS+f1syRHki7A/EfMXAZHPVTNdUtliJcrOnqs6gJ2Rvlw3yczaXXD7Cjq6iMaR+MR4
RPzPd6MKa/cNwwH6XcZgb++7SfmOIDPyg6GKtGPw5t4M9RWt3tRFdFbtpQlfLNgzMQBCLJzL9Pre
Zu1+wEL2Eci6I7ruAJY1vnmRokULJ1f6wv14FNiSVB4rBnsHNB2LobFauE5u3z+ROcJD+bLVMkC+
0B0zo1YakTTU7cab4RJVtUFV/nFSVO40lGixaZ9LiepYPVOSG5yXI1k0HaIDgn0ZK3Xwf6yU1clB
6gSMVUoyYDuuCLI9A8vwBf2s3W056K/QzGCt5m3Z0WUuwYwTlT5zayZSvKCqoiRe+6uL/AQkZ02I
hG67XTyCipaqccOgDVbJEeXXP2tOC910+W9J/QDXg+/Zn1P9265bfXGJACiSsPL+GcjAA5zBZ1NR
ouTKI0bK8uEVlRVtKkUp7kLN+ncnvQ1GE5O8a/71bj8JBh9EqIMO1aV9K7IrUGkrzwklkJ0iXjZw
CFTh2ZfziUrd+oWSrtjbNR9fLGYe4J4XwakiAso9nkAfVJMkQt9kEk1RiCr1ULBjHmg9K47yanUR
RhLg8aIO5rDMWkhKN13J7cHL7RZkx+GwdleLAbiia5Y2cj4dSur/ZaXp7Vah+i8qX0AxFczQGhqB
C+KLmzqTaaeGCpTvHlnwG2ShR3VCtYdRzMnQeIrCHTP+iSADtpSG0ru8NhDfqyXI3myWFv+CH2lL
uPnzvEU6QKyy0wbdpax7iwxWV3eL0mtzs6Kpn6hU3SKyANpPmaQHf820H0c1ELubkfyd0/ChiTnz
TJDUsC30FLsXoGQ5tzHbftG29njClfQZ+cvN5I4oJ3ElQXKLTHhSmuTCq/9RMV4Z0jt2PMk349Ck
/gV9WrR7MAgLXlW/YfWG56UMC6bFYFrN5yqT5pjWG30QDdVGD9O0wKFKoJ698wG2AOS3wF9SMQm+
je3xcIoxdSOresYmzHjQL1+ZONOND/IdwI+8O/OEfG9NsfHNuoybDjAPW2CJ7AJBliMxWjW39kbd
EwZh/23d3PAe9EemIOK1e5wJqRu26b8FaTfkRNjfccNIv4H55BgFey9xBZXAI9y/pedCXOai5pOo
+MbGSVVXwR5lwSPIiClbglQatVyEb7xItL119gBe+RHnFa9pc8bvY/G1Wb+il4Qsv2JbDTCTV0cP
HZOBGWLObmZ0jhPVNEKVd5adkd4Ij/ZHFuY/2IDQSUtndxk20SHcM8yepyk1Ko84M5/lh02z90Q1
PZxHIHMDnccH+wxmxijfnn+VIyIgGQF+0r40oQBOSKsstMGKUPTguS3EKQi1E0cBWo397YiTZ8Wx
/JRidTfpezNQKs5JEtr8Lh3SWhwoSKeJ60+0Yg9Tr+z0ZAkKCbt4rZB8NJ6r9bspXfJUc642sL7E
J4x610dLB8OKdOwwTWpaDE8z3MK1V+AmKasSRWL6Lipu12GNzTt18W+/OINAxerTJ1v48MU84Xrq
RCvRoUxM1MisGkEfY2eiLQ5e+UCFy5rvth1cim5py8/5yU6p7X/OvLxY2eUKcBA7c05SQiN+O0yd
cn3ACn8XmpPDKi1ZtodIkR3kq+SgsARWIBMxndoFfN3Q+H6YUnN9a1kFXZWZZebD9/LvA+8N5YL5
/KlRdmstuViwY4suJQhQ6TGe+DO87Qlo/qYYb2ORqNFpwZs8GLlRZ4ONLiRlxn3e95BjXFqrnk8z
f9SnBhWedQL6Oa8Lh9FjL8oq0+daSqP+mZsgbw97NUVcAQPWLztnU27wj+Ez4+EoaX/V1Lm2VQSA
IsRiYFaEZRhrX9C5mDFedcnBFl4+nEnJ99UxpCkHSTYAYTsfs+gPkLnt9BKvv9y812UVK75uYly/
zCoP69F1B7qxzEw0i/Ruy2edE8jbjMEuIQHjXYuoM3MjSrZ+Ks20MQPeecJkX6Ml4NugPPqFpR85
2cZ4vdrzfgynu3WoJjBTh1L2tO1ksLsHnryp4lXXrpXsPtqssUQAqWcijxDYUuSNK4a0vGmnHD/+
EsrpNQ2Jw5QZjzlWnVXgAQERIFSPz8236eWyMDpo0N3UsQmJoZmox3soqzJh7gwF8LIb9vpuZCfd
/YPtEncQXIESc8bQPopUcTdk++qkTfzjZduYG6liotex6Zf0O6/CK/uJCjdYQIEd0tCeEsDXfIuD
CO9LZx91LEf6StyNKir5FPD/5vK/C/I9/6lEOWaMn1myPkyX+mCti4kRlsKhKibfKZywjF3gQM/s
d1+KQu+C/OMsUIwZQCPMV8WX5sWfl61YDZB7TWbk8A4hhEHCKfUax8dlP1XMsdFeugr8lELd3k6A
DZuWiuhb9IzSCbw+qmlF5he53RedV3GNuxw3MLzxuuV8qAsMZDnpSB1/qbc389K8ypsgBKL0yJSt
13hb37aHbwtwQip89p6fKyraJnm6y2gj0awiYT++cefzK+xyKLmqdtT2p2Y366oczQGceZemFrQR
tFlyTdq1J3naxmnT9b1p8NGbyr5bY4yCI/5c8esnsa3jShB+WGNM0yy1tH2clqQ1h0XgjFSAZUXe
ZjFU8MGkMJBBtyfHSGpbnaKJkqR7TWMjOapn3GUPwFhzabxL/h/qAXqXqsOv2GTqBLcNTOtmAbbv
uj9klXxa0Hoe+wZbnoizwot8OqvV4osP5QvrEdKo1cNQ0W/q21iKh+Kws9wCAXz96p6nyUsw5IoI
/ZhJAGlPjCHmnnd5FLGjQD8Q3Txzk/nLy+g27ZbarANNlU/RWH9ueilFIwzMEjNC1qoXmEdoCOMv
vdagSN91uEAdN6sVDpmrckNr+hHjmWN1g7aZjx1Ps7XNw0cXoNQmrGeSmKeXlEDKFGlv4w7tH712
nVtK6gaT88XTfPIjuMuNoDBoH9KIIiVZw7Wje5rGy1wScW8AU9cmqzwnl5MYpiX+WULJNWRCS1Og
bWhN7UDzlh0kXcMkXn5CuvDHR6J9KmxH1CF1MFJly38jjQ6lJ4A7aaHg3c/VYBGa4bGDM/jh8R/4
XB2poNoOYHiHCf30jn4P5JV1whIPboYcXL379WK6fI9YnFHk7rQ4JnTssx117hLeceK+q8gZ584d
es7RAvxpx4H/8F3/wmYtO5ib49zl292A1CGl7o+dpOXlGZzcwl2NearNQwxysYbHd49b8QlYUJNh
bUFZsmpjx82WyckBL/nEVa8UEWh9xIVGv2wX1ZEvLNDcLr3xSCr1LCnxb/9h2vM3ZTsBOUl/GduX
zXP4Y7CEDX7Znsp1ydQ5sQ56KX/iECitMLRVPQ9ASSi5LpyHM0XYAXVXofaDAGHJv4Z66X75EhS/
q01ME9OlcofrB8E7vlj0kdZeRHnaoZORI1gDl82E75e7eq8gqI2ihbrIf+Ec0luhMTwM3uxj6seH
w3eYbUF7jFQo3zIuh/+Llg6cEaTVd54Kqsc3iLIaLrDaJcap1AB1j0Zm2/K11yVRfFWnkjZKAuN7
ayUMS68J6+wFtoIWQ7/mFqpjpPU3pUBS65BhoFmEGjyDgAHkjmOxUXhb4NjznSmnzqnTVu/M+msd
yA2Q3IbQTiwSpPwjYMM4Mo7iM/up55F07gL8q9Kaa2oSpK9l313uDuaWqYvdlWtcc5ht/eYwr3K7
AYTUqBUMkufmthkW0FKEBmK4/FkrvDS+DCV3kbgwUES1XG1DAVM8O9wdM6O/88AMsHiZYqRJ5ir0
8+CRdO/+2T5+0D+34n58kylzfTNXks9YYsfPG+KmO2dlUljeAVnZE9mUMplS5Ro61UwzLa8MsLjV
MBtnDicO2wm0fFPKGgCgH9vO6tnjDg2J1Ysz2dsDIqNcTFWyg85R7037gBTuew6FTaixxwZpjEjk
OGbbdPtP/l+d+Ml3y8OXdM9jvX9lHYrKNnkkyKJdGFIGCa8RW0IubEc0AVUYLMLT+B4qOEPdcrc9
u3sbz+YNG+mhCKgsz7hTZAqRaBEKH/GUQxKOhZ67Ujd+6kAP3oVEtFE4xuImMlIGAYd6X9cVP8aV
8fnpK5mbmhZkxS63wanG9Gwrgnycyob1d3AjNwMU139S8tzBbixTKr4l+gf1VqhimuOpgloRCqmS
8+cAsy4k+zGjeldFu0u9ejNvpak6ZgqOUORS9g9toa4BDK48mhUFew83r+GG7VjeMjv2UqVcZCZa
r0vKT9dSjTS4Wg0Pfh70yi5OtAXHSLGoY+kXovG3gaUCodKACfuPUisx5dUZX0fp8h6Ujn/NZPjv
CodSYGaDcW6lWWM+j4Im5bCdAxF3yaTvVKccUZfnzUFYi6gnJpFk94cQst5nfv7UU03b4F2m8Esw
h2wb+BcdM65bdzxu3o6ou6z24PwGwR9FfSIwmL0FSm4fAOx6WGPVYszzl6IAMDN8CosZPr153okH
deGGbVZ47jn8+YabD6T8rm7xLP+/zv55rPvIArqcYElE+annZl74lId9y3VIl8huV/DaICpRU3JC
QAKIMucwct4xWtS6jt8ypC509QaHMaZlOpKWVDCoc7jh+V0HsXFbG+GKFYFe/NvkL39NUTKXQw6C
Zf6Z02AsNHWmOgxRUMqSTS8otRSxsoIGE5VCSYmvKhe1lm5rRvShJHHNXilg6D2veFuRemd7DBim
4YoJLWcF5db5RkOh6lq4WAT/CkwFqkMx/IB28umn4ViKr79j/QxXOdMzP48RwNH6g/tyKs+dO9Z0
mVX+CLBiCbLrk2Pd9T24jT7zxTdcD3H5xUDPqQQ21ffzVUVnYDPIJV0WLTmAU1NgN/jngnCAZdh5
7hIl1MWBj/DTe9IxBRIAh+P5AZJSA4/2QrqHw+drPoJ+6O+pOBw73EiQU/pUJHiJAlk7LhI/NjtB
a3m/1K7/kRoVUftryqe/p61yN/UgMPHmZUY5+EvoFC4RBBd0NvDtFTXAtKI4oUEoz4crHZePidJe
EUPwHJYFs8ZIiKEZx9NE7D6Me6rPBbMcN+byBngSZ5ETSNFmOSi6wm95DvNwAb1A0Yx+1X/s+Yur
SZ71ALmvz1U0bcp0uRsaHzA3zJVNITcBsFB9T3km9VJVZrMDgtHFdfMrsjHfT4OVt5ZjqKx9uz3/
Vmohl9Zdw/aNWtPQ9XBzvvAR8TtIJLVxS8EsQHwEz7mpYaCgRwhm3722V7ajH6ZXSe0iPXnzbTdH
9krSGTAptLJ2/MHKpS7aeXKxQH7LxlAMIRDTMeQSNeoF11VuJDxB8nmq8z1lc7+GThi4ssg0NdtA
W0Ndu7jelXxzmgmEu4gOJx5og27vZCyLPmZMaubCFzJQaYvnYBDMy36D3wj6Zp+f/47ql23Q3laH
bh+b6Kux3q3siMATx7C4Qnerd9pHb72j9IUyPQigtO7XXl5U85cqbVNVgjWs7/DcYMh9s1+/Koo9
RB6ebJ7Kf8IOSsrd9JZMK1J3+dL/PuMkjAOcKy0R/PzyGmqm0j8cjz36IzgXTzcLxSZKcjmvCcFK
7trU/iB95XO6i7+UNYjkOpSc2ej3kl4pQVER4zJFLYwwQD8y47sUN8A90rSzdxjpJF4X0WRRPUy+
7O1xqTf+d0rIYzMCLzcxb7ccadapxBCAegtmV5jTKpZxtqqlulDzhe7jGbCcvDEOXaNfg3vs+eF6
41U5Y2IkEfxTxfQDRXVtRnf8L0YZNTAEntRXh4aJxp7Axxil2cu2y+Nl8r7Fr5JydBpFAMQrMgY/
6UsxU46yLthXRh6FDvr0q4YgR666WWZ6HQ4fxoIxc0iuNCCaaHeSLMC7UtE8QfS9QlAfdF72YYu8
CzPglXIGUDFDH8KoBJKL3Bkd50MjI5cyJLhSQSNHxK6T/MsL/FLwjPmnYHjB0n9fRc1pZNSNarV/
6fJTBGSVMV/solusjTJw1NRlz7rEEHmIJgGWO7c5eyL+v5WXY6eedKU/LhL9z9/FX+un7T4ckh/w
NIZOJfo7HiRZkfinf4bHtOLuRJK3Id9rKTJNykYIOLqdFXiaG11htx4CsEt4gn1iCVTGS7qsLsIW
tJGD4SKwCU37nWNj7JB+joAKisGAGWOCKuwfzAAULccNDBgWcWfbxfL/ag49NEEK+KW1uXDaPSCv
7sGThSdHtaL7dB8b1wOP5DWtt1/UOFVqlrgKZYjvAJnRrrZxpGRFMQ1C7DPkFAShKV0lrpt1G0q1
boGYhi6nT8rkVo6Pz8dnuytGTYYcmTGcUamURwsWacJ4ZWQ+FzdQBMC/lr+0zBVf5LbSjSHwb9VN
3D8G8kPPJhyA1009TJA1LCqezut3h3mR2jEG9MLwEhMu0i7m5bxbhudZeh/pCMBL/hlS7EjEOwkf
mtTe/TT8lJTB++isl8t85ech6h/ZkC4Yqp+hOxBh6tBnymI/LBZZq7Q//3QTUk79cU7SGbJcNddW
ayYFOm7u0+NKylxuFo0DKGatPyQiqSL/lvK/TnetIpHqKW6N7G81Rv8udtdxf784fv3sabx5efNv
tYHNI58lSVVQFx/9pKibN2THmIHRxMjoIOLlMVStpri/Z24X7N9ByNdYn+mOjwhg9Gyj/fAi8cfX
hfNQF5EXl0mFpGebHYa+ulHJ2qTQFB6q9Wjetc/gpjXVB5KrHwYJbFA9lyPTaQkrktyioZMFyH+S
fwoZETLQJH1RStULr2FbGZMrLCCR7OM/iC5go8qLhtjnB61gVbCaTlEqWJwNJwvqiu55ZPQdHYGH
swaJ7tlvfQITARMputih6bWn4FDfJqleTW61hDUShp1kB+m9YPPU/KhbyFPZSzlG1PhuIzVmqFk5
Rj4XcGs5IiUlDzCbMlzbsT/jQ5irhg2JEXemoEvkh3kq/WdVnHy7lLL91FZPWbvaAW7oek9nWGTZ
sZOqdyUQPLTc8dDpYmKQoFTAvbGCJ3+DmZitR75t6M6ia6J4D3zztQZPt6vW+RvdIshNT6WQO3pa
Da7H/iFRne295oYWKYwXWspe7EY4eFN9xqp0vwZ6Fpb6U4lhQRcxfY3+H2NFu9VxJSzRlGozkEsQ
QG6F4k0TT6ygUtpWpTNPWzJAgLLbpsSXbJbSOlOo1CBFWdZ6wsr3txCig3uJ1mhvqoQwABGhgjYg
p+7eoJk5rl3n770k+Uj3KZFzGRCsJlgl0YKdZIaZ8qqlUxt/ZliIi5jt8IKKX+cz4m3EjwBTln2y
foXob8N/nHM6nzTYBtIC2TOdS3UnNUrcY/sgXVfeUuzFaBXotBNd/PL10b8yap66emLUBMqb/brB
3nepFf0EaHXU/V3JsI7kRVdjZMYG/V8NwkRvNZrQ9xQ+0iTQVaWk7YRe3uuRHg8UBVEGSDB/iGG4
0m+Z5LqadtG/RrFL0BIxaOczfiyYWDype9zTVXoJphP6LPsspX2Y+hkxFu9mAoAbQvcRr6a58wwr
G/9GBOYWOKTO5SUUmMK3CUghdpJjFZ8kpjpyrQnGWCvPa8h2V0NIu8S8ajItadSi5sXLwiCOK7GF
m5nBcWv4HJZmbRLi/An78pjmhqvRLASlBQUwWobVhJafLpCPeeiuWlMoo0sbAlH7Fj4MRemFfG/x
qbgMmjzHbYr7Ws36HXgRJPo8Cnb6y0H36Zc7293DyzhlnN5OMmfWfxdZqc2bPr2oZLO8M6hopVxk
EsOUCf5F4w9CPZlmUkmLBhHV4Y+HnMkKpwVOA1md5Hcnh8g8jz88jn83C2AwZh/OHXfSDBgP6rkU
ZPukylG9ZZeSOLRZTbd9mFuWLkwsWV8t8Y+9flUXeyeNWSh/hQsf7WBCOsMswOqJeXACY/vzKLb2
c9eitj0Pqr4LWNqCr2l5Aw/3i1UUBZWkNSnsskEpnscye3ok8FgBegKeyNpjOV7luSWV4OW87sWI
irs8sGuvrBVjSqWkX8AB1ViW6i2y43Pr17l12JKj0lJQ9jSr7eTSZzymgKygG3lFbzfulRV0DJIA
eJF5Z2g59/BZFzJwbFNiPdCPo29eb5ORSpOxMRvdVFnRNMPPHdkJrk7Hxm3k3PuulP4Y5RQFezF7
hZAWnq4mNPR4Dqu7qopI9Yo5PByxSlYo2uoLcuKLwG+qjId+9HZI9PDaCFKRMQg/DVfG2ANzgWIx
l8Kpwc1NKg+o8USSIWmNOwGKKauWfXjlWhaYt0APxZZn6So+OJLNtqel2Pa1jkU8ZUXTAlmIYwhV
g3Rh0WKE669wTGKxFq/ifRM3fxy5K0Hl8bT2whz0Tpqfo0Z6mGeJt8q2vZY9dx5bYxHQXKaiX4TW
CqMX1VUvdNenc5lVn0iAfyJcCBoDybH0AQKTnLW5G7bbN/1LhNXntxAWl9mXTE/Gd4S2ydq7jRVG
9Hfqyl3/PhdPNMQ3P8Gq+MoiVlS5o0pPB30p5AQfD7rOEg4LiWpxgJJHz52EhJsdfLQDGq6Twjhn
RFSABB8VRoBRyfWaAftLa62ydIKfaSrudLTEeKypLqTm716Dja7osUSBYKl5+dBNwlUxTxCH2vM0
j38At7ekbxHyvB+FnsetXC47CnXDqlM+a2YIami0iijRg4Ld890PW7X1nKyQCKLgpv7YFeAbx4Lj
+nzkrdlbFo+0DSde4waO8Yhirq1DYTiXnJkBzkntoXWraK8K2deU5wHj2Q57NrFxu58+aE0glPIA
bzlDdU1y6Lhce8IyhQvT8RE5tYFWMwb9riNlk4joryfoX8ciJ1GNabQUJYwBFVJjLbPR25W/Wb+B
WboZAgoi6ycaGAzO/WqGzg9nEcSXQ0ns43mjeOKqgi0KMgU4ZxB4ZY+O/oGhu4PXLzKZL7uVeqqw
Jlo6XzX6Bn6Gfa+AL53Mp0B2YIedvLKxUwfae6vspr3nDd/rgL9m/8YJoC0S1ClXg7M+9USjoOfq
yATFlFudx+JNaKwLSafwy2u2pFhZx2Fa/XCct5ldzi+B6leZmKzUBwlerfHAjYBQ0nqQCIOtq0Qs
aoR6DMqFHuIOGtGQHcx2IPoda2TNoFcEeGH/t946TqjATxTCI6jyQtLuGuRlKpWGewtlzhTR+7/T
DaVtW0e8ChMiwkTWWxaoB447buSVtDVeiFZPD/eev8Y0Tc0I+u4th/8fQi1hYEkm/ZImqC4DGMzA
tXE/2RyhlXhnhS9dVUl4hecwqsgtri2Q5LSrAVVwLW+jYnobuTq/ARLQxg4Ylqlb+1o8KtlAtwL0
PjPc6LzWWbKkUpGLYj0A4jN1VkTbDQUuzUFol1hh9jMM1iZgWznEfexwOTL5v1+KJpkufCW4oL2u
bwE9NwokxV+jJb170zc/4n2B1F4pLZxRe7q4uV5yX26XVniA6GpdMt+DVEZ2AWmDY6QkW1x+vnTb
FG4QQdzRTEuHL6oAJWlmqWZ0o3Id8hYnez/8jZR0+W5cCGU9Fowaf3cELFfFYWRmV0SjD2c6CAuK
sqYx9Gp9S66B6boddStG7IJD8eq2A7H8wMW5XXmQWlVSEj7Mney6mSIAVEPsU4CchfIWNq0ud5W0
bKn6aAudBF99IeNNB9JDzHnuo0U+Csoi9d+HIGIooVZpoqbB7FsC8FJ7REowCOC7v5h6MFNQQ847
d8u3RkSBExOVWwyyWl6sM6GSpRU/mAECWMsy03AWJKh2RyWI5JHAwReFF8jaik2djg+j89jRN39f
03rS1ekF0mApoZ9y44OVKfREleMaJHml07wT9B0R6Xa8n7qBQnktOvlOogW6JKR1gV+bOZqHvQxI
IST2co6nBhSjfkgK3vE9M6wK5wLuY2D6VLEU20d4YCLaO5keePZUhosSV/SOFB0Wmb0HA/eFMea9
DgEus9xJY/Y8HjZvGDHLS39WrW4BLNeeCJoO49fWc7/Qg1Fnwju50/dkNXffT3sg99znfIQRTPKN
6qebBNXDGDodmtrTo+LHmdhRJ9SAaKQIbBpZZzKrRB33GiwxEu4mOX9VbQWbt//SbaGi0erCvEUO
V26k08I06nOBXK075g2QWJR9Qr5wih9c8YZMR0JFUov/iWUZSmv273WQI08nCLK8FxAkdlLU2T/P
qucJs9OvpxMxvnf941kOafIXjtJ+7HLyTTcgSFudkX3S50mXw5To8p8l0OQmLIFTWxToROndUq66
LNspzdynjFEucVsipZjw2Ed8Zp1mStFSuA8Id4K31y9e9Jh1j55Y0n6kP8r2msdhpFHLfyVzuRRi
XUYd7poSqg2P/sp6eGxEAT+JeNve2rQDFxv5NmyBR8rz+vtfVhjkMvsQLqEn/H8f1HD2IKHvv12O
duKJLzGejopMRmhqwo3/fR8bBsicVuLxrAIjgOCJT+Hf3IU+pZ/t3fg3iDDpJMax5uzqEyPr2obx
L5vd3FMI0dib8UDqMVDm2o/jaq4bRaIFQ7CnXKW4kkjHToXNp3yxLQe5iK8t186TeJs2bfh7bwjK
EAWV+rnMlgeMp+jTtY7rUiIYYqM4lneYw3h334p7DFWUi1T9Mc6dPL5jr55QElvWCKyIjvg1CrQS
4kRkjUt4xwbw9Rpk2Q2NMu4uVOCRHUQFipFCptu8tzbxUQHcPa/JfG2x9NEqWdF3saqCfCMrlG51
IBJpHMP5/Q578KfQo2AifcFT3RM7jpEBJ7OI9WMs7gHth9VR0XJ+ofgmhVHY5jfscwGg3apxZ7ER
WnzGdgdpmTkhnleLPAqb+SLsJJ1YKqMoiX5LKYnrOxQnTsv4E7GsSJwYhH6N2kXFpSbI3ayfwAob
luw6GPeThKyYKlwP9u8QAfpIxl8/scOgeqtmypObrq2Zr3l6JXSH25DIwfOFh2NODaqYqpxeG5HF
HZsGXRVUpmN0vNCTEcs1PS7yIkKRCjxMU+W8cDQFKyqsnFaSM0/9+x4hViL7BwsWpqBL3KcJxCaH
cIZjfeuEKGIhlL7/1prSxJNxyyepnooMIsStTCuBECcbZN4CqGYF6li3ywNX6j/doFHW01zd4arr
xHfvE4o/4Mwp1xHGdcogI+imbo+ltY1bJVLT0NZ48yWYUKWFnDpoa/E1H5s+L/j9xW8msmfEcRIU
WWo5kGcNYpXvBGfGWiTf89xCVwEXa1MJxSZAp3XH4DI05UrMwGEo79Vv+yYjbw14SNVJpv3NtKNj
/I2qOVXkwIUzaZiNrHo4/Hlqjetgra+2nkzVBrGpL8f+P//YQEoP0LeUmIFP8P3QZ6mIbpNaMC9x
o2+Ywrkl+0skcKIT9nLGxc3JVnJtXDc+NjZ6xemkv/zPQwb/ZHAxg2eTKt+y/CF7LI9qfaUVibCe
RELiSGi/gTc4lfnIEdZdA2l33bbS6MdYxFO+sQgYM+GI/GvcYPQUXYOp3Cf4bBriX80IWJhgAGqm
nUWNl6Q3aaoRuwM7u9UJpxJQpFsV52vQKRDLA9h/FE31EaTTSiXMiifs6s8ejDtAJ8/PZsxaTrw4
QiCHslBYi2fTflpd8gqxHp96mTjrGD4Ztp7Jlpv65LLVrZR9BxBMB9u1S0vo5bW97cx/YYWJ6nvh
92Z3uimrTmgyB+wtzfBdZ5xFhK4d9HdiOFC8Bdy91JVPri95ZXoidISo5YHLlne9nsm7JXGOu3tk
QJjqarU/7qrldfa0xJrPwUkpmacC9ZTRZrGimO9ilCv/XsDRnC8LpptLRUvtkqRnTsDW1+31971I
4PD+rWqOyZWDJxQKfStw+5eHn20bjF+cDURulM9gBceRLFbGvmyyvdZUtnPZAkh5mshfb8QzTnmX
D9WpO7vQWde8SuithIrW5ut3+KeQdUBjw0pGRG/lr6hDheezqF8GQvYDX7v/EGLDBsmJ9gCtQX1q
jP1f+KuGqlfXFgc/GWw9Wo7hhf76UJ3/C4Q9qcgyxj1tN2iGfFqrPSG1pwSNxinwygY0d57S6BpN
SxcA/dN8MwjgLCpfWU03AP7x+XwGj4bn573bXteQpBH/BJE0sixez8ACF2JaYlukzVCv5YRTyfq7
REMzx+hMFyZcgoKomXNyt7odZSlJmGlacgDxH2aCJRZy4gLmrknUlt4lAhVhYuD8zX4bEKH3QGIo
ULw1guc7QY82dboMWU+dudmThHfUoJjWteYQMcK1ICdLOK04g5kHz36QKRKLOyH8qbNhFdztXMJh
g4i4J8w46ir3c/H/5aIyme/QAHiXcphHulEvaCxnCMdC/UzUcRLZ73sJIHiJFzQGu4ALNXx/v8GM
udZtDVjGvgBUyVHRbwjAd6l1hYR/EevhZYXyVOdfBMU4WiOV12AbYJ8RlDNEow+mIq3uqx4GVPmm
bvkYzn8mYItne9pVtEECXkJTOa+sNjO7wOMpCfBNUnxxQ8L/csR9ZzNISfzjnTUrdg/IdAHhWJvY
84GuoO+xwg1auTh0E3e9Gmy2rYkw+5DugMRjfvVNHZari0PzoLSVOdbNGpsfq/blF2PCNwfJL2Rh
52OyuTsbr5TXPGf/V7Y2RcK/JbdJltKF6KdcJKzrdRUIZ6IweV/EtxJvFbEqZ1xs4bqMjwtyNSAB
Pmfp84qoGBZgOIKuiQa+Lquy3C7Z1OV0Sl78/nJ3ecU3chAsEWRkB65PClTIRxVW7SMVyDCCUttl
bCqNPSxAFK66B3P5R5BkPWQa3veza8b72JjgOkslyDB7DdQ5fjyD8UFYIzHPamu9ucHKoGcq5sCh
arzINzJYvLCqoDwi9mA7gSTUB5UQQVVqL+DOokIGg4Gex+b5AX78rCF2RS13n5QCJH8ZSENoh7Vk
jxmPrjHn+aUrWBMpB0NkEBqJGIf0Puw+wYBHZjZbU9YqI8QZRVX06lqCkQfPj/zahcWlZp2Yjyuj
2qVPlwVJh0nv0nBZzDD9qz30rjm5o0QTdcPolmiXF4aan4wLqlCvJoPPMDvbYBS4Ug50bn9SSlQ6
gKbub7kBWwemJN8SQMZCTaQeuy1XK5RGOqPPgIoD58BRXrGgpPMu4erm67scUNbW6gvFCtc77jrX
cW36O+wN4os1kgRU1lolKHcJHrH2DyoOOlASoZS99FgOI2puJNx5HQeuxtI0hc8ZrAbK20OkpNuw
1vuACNyc5M9QKYp60ZlC0Dk7SCZEVkpwJKxpz5vTGEvzfPnoAUorU90Xfe51MC7wOepFeg8goILg
doH5g3iomkNtgTSxg0TgoIa9laWYewbxxQ52VIo5FbPJT24eXI+aSHtuU7Dg7HubY6UQTfDwHCSk
jfmRB/y8v79d72kH5OaJKxOZEmelCuWvfAPGv5YTz0Vr7AY4Jcr8cnElLByUe3RmPzhN71urG+Ot
04mqkl8Q6REDS9u2meHH4SGOLxUHUm6r54S7sNDAAlrRpp+cjrE03Ct2IxCGncWrj4TRMU9e1fcK
FvwSiqOdvl3UudWFJrs8PrWP2ATYpQmgnrhCxUcMHZ68gak+1kjXZ43FcCbzYr0TMLFupqn88KGf
KQwFoupzUux5lqRAUHaSj6hlLZH7UVna9HcPlqgJ9y146/ebKn+FuFp30OuDqMsZ7bJVVJEJviVx
3T/J8+owVC7R0km3OuT4o5H0E2AfeM5HQUinVJtvGhlWYEUtQP2GZ+Yq63TwN3PhzoyZ/LE7PlBl
DX1K8D126E+yc1/meeiEZELjIXrw1cbjU0bbrMDmBep7tc3laFnuSQ9kz+IRba2O04udQZ/6+7UO
vvwtTa2egoPw7hFtEDT/8rCvY0J1dqlsEu1Xl2x+AHOQEU6lFE9rwQxXQxblU/WSGW5IJz3ZOif1
vN9CtU+9Diy+ByF3ssDrnvOa3emT3HRnX+HfI+wLbGHoGrndLEmuHJNgnLIhv5bI9EXJf+LKstnB
MjlOcyW4RUCgOqcZbTX/XfJcuR2/+UW9rxx2Fq8d1RS1jN6MZ3s/m8XsHzUxyZlUHWq7BcS402BN
2FCh1HhKz6wRy5Sy/XuSvnRPmoEg2eyx2J/1FmMnVsDSsxlxH8ZUBYhOOJMKiJ/xOIoNM0qeWhyt
TCf3BqCCpFriraVnwj62+A4JUdyazLSE4DbRNaUgtAWMtgEsc/5Wc9/YmkWfvkorzeXQUjJo7Az/
ir3W0akWvyeKtxVk5TTzIuwy/HUo8rghi27qfHm6jZwfns1PlOuojjyT4emOJpcQad7sqi5NTI3/
wAvUqGxF7We64pKhtlAPHpoYGYNqP3z3iuTNceqv9pTiRvCmn87p5T+1qYOnHyK6zXPd/TjAp6rC
t0rVYyNKD++eflT7YgPNQR2EysYGmYSGSfehNwxW/Jiga2ZG9Aqn0Ya9ZkjnqTOoifhEur+Or1xa
pDwcLKyIYFv3p/DurBye8ztjkW1I1P5HjCUipeEgepq/4gR9hGppvm6qpCDs1ucEYzh58XGYxFtr
9+EBb6UaOuGzfWZwSNg0p4/8QIMXARcqvpot0+CmyNdi7joL6iiui5GhmzbI2yE4eyVg5UU2CgbT
pHmzSVk8qi4InN+noqVuPRF7QjEkSvIhwNq2mCCMahxX2fPqptd5J8rFeF3iBtz08vldPhXFzsAZ
Er/cAvn7YPqTGAD6BAtPUcEQz/NvS1V6Ju6NQdOvBq0ppao0CHVtz/WQmK58B6LMEjTXV6FA3qjZ
7ykQQJxqsdT35M2BXAS8FbmyhK1kf1/JE2OC7H295bXTDqABRdjtwN5vTunN65MYvGHluOeDdIc6
uFHpMidwlAfiTsqRnL+nta7ZLGuuKxKDj0LbYMeYcDs3Ubsmhww/sbER3aEJsw3b6wP9wJAKiySs
4MGRg0bdWdd/4zHoIRXfQRCB0342BANguwBz9sjEASCWELGjjV50n6bw18ov0NmisEKgbSCGU/b2
tPFj+5Zk6yFm8fez+Eyp2vY9xhwyiSoXUOuCwDiUgWNjGqkAuibF/pdilQC2rWtvOerv6gU6IYb9
YctK6bF5AfA4W2/JVT/O5iQf7Ku+aIroJUGMTRlJoerG9mixPanSxEqjQHvhgIAt2v7jDJv8Mgks
tTLxf/rnNJbfne59yEj5gfXA/9NhbU6Tzqo2JOeOkoDmxF+9glCA5V18w1U1vbzytpOBz1SpyPz4
U587d5LfZ6P8vAKxluab57Hs+KNDEGPpC315ecLO2zZHZeVIA7rogU6MHRGgff469xYA8I37k5I9
JX9XASzdMeIpxE3qhjN0hScCZyZtD4wZBO6ZBkLIZewW1rB8jAHDV1/EjAFZ+Xxd5/1L7nJVaYVq
tToc0/zWlEX667V2u5GPFYurmgJCpyMKFIK6S3Ay/9xt9tXrndR+lM+95N+i7ug9VZA2fsHQqBzJ
6fo+v+WRw9AwPXrvoVEXj+r8DqLyp0+lCv7lBV4Qat0fbWXHVZ9x5TxM6MNjk3TSKwYIb9+bbIW3
VfH5QDI6krgk5gTr8gEru2s1tTzRAU44ag4TW71jOoAtlBNbauu925kL8x8DBpNoBKBfDug7Qf9O
iDm58XNRPq+bvwhT0bPNRCwjy+H8kZgudHJz9XAj1qBJUXLRUWYRLgEWqXxmFUi6HwkV9IsUlTYL
oT4TdYqXqOapewzKtB+il8mFNF62lomztZuBbybyE1k68Z2ZZOzru3lwBywl8GShMOxYER6QQaOn
VMfEoUhj9oLx9JmeOeoHGzr+eWoBhAgXZeRCXtZP7F9eTwVvQwcDuhqJNtCHRZEY+CWRRyXZFcsz
Fbik14qOdQib7bo9ISOEoajO6l3wQBbC7xPqkY61SeIpgbjpxipDqaN35kXrTUh2Hku4Uv/G0TVR
s3rNS1rOUAmvz603aFz+q/gOvRi/hwz49o3Qb5a5+uLA9fnMrwVVejOHf4MQ2CtwBUACcLKcqooD
VcGXO9RbnOCE4K4tItUR45nyxEKKDmq0F5+hHGwC5XD5DIukpJvK+GosYr5Nv2baALKUrm8uIynF
29FaSPS0VRe59va53QcKv8HeBHA29bJmVqLxCSujSorJaZAfwvNRt71L7jawqgUoCSWhiLsFpyvD
1MgaCqKeiPa4f2NE843icjw9UUE9EnXwjrk5BPyJJIZ959YzRjXI9wy5apHwBYQ+mGRHqaiLnhK6
D9K3+ESvMxoWbDG/COn7BGeDMV+sASAbP4LhfMS8Rxju73vfSs7C089unHytr4FNhAoWdbmFXvVg
POorg17Q6pYj5uXASNc5/t06KGnC1E1wLTni202G1l8LxXuSf4wEKnDEylIGZRBJZIi5tYqROVRK
MZUlFC+GQUyq6Qwohq1+MeDhsEtvUIhvxKOlBnlahNIRFQ2PCkJQJvJOteNALYdejzhneTRx5RQ+
dMprz02Ui0QvzVkyna3PfHNsEmVuN4T1hq0BtBTHZLxVD24XyNF5jUy7VqZt/GlyrwRsSD/IU8b7
1xSOPgkRtuu26hP6T1mrcSyLRdgARwVOZeiJFWuvCe0EkE8h7s2K3DFGV19dnsEtrqPXAgRmVOO9
ykdtQpNFdvwRWWT+51jlHyWA/w/eKPMmCOIl5IUHH8vxPRjU+5mSc4kUcTj0G+nafdmUf5iVV+km
nCH4afdaT2Gd6KzEAreGBLF3zTUciPlzNGfExwchRacrLn9Mtst0APr98UwtbsUtYXgRDODOrAWX
vmAp7uVKGQbhLEIN27g5XgHjLQJDIgcvRYlWTziYduj3J1lWC/NPpKQmcqGjslvWEODAOIVGEm9A
TApB9Tc6YEw5obO6XRe18RIwquY4M59uZSrk0HyrGC5juHcquQLoHyjltOO4PriAc4lSn0oxkSFt
632cy+JEiDP88EbbNB1BZ/eH1bDl+tWdwLi+I4afAErAx4dbHa7kTVsFeLSnH4Rbk7fy7fMNcBqC
Vu38UUEZEPy8h3x8iAAzjH9d/XyYvYYm0TaIZOpIPQ0u2uZa7Q5eHmSQbwSqqQmoVRchjEsGsiii
FAh3Qr4frk1tCV3lSFHiRqWjp0dyOTVtiugZe8YaUlQD796jMtGhc5q6uCkfqjVxH6kSCPZMIqLF
7nwRnge0zxJHiXACCyzwM6vhZiO0iaI0JGc3gQfpnD9SV2C44K2WpHW9Jd0/U62s0LHjo3MvviHx
cfUHXpMN20wMauZ98dVwaC2Hvkvjq63gWddUieAvHWWE4i6AXgQppG+bhjtzZ8gy7icodBruex9F
gfjtLVp3Yk6WW2Xsg/1jeYWRS2E0fWmqdHxsoI9anYjie9qbk4G+4MPqlAHDUTFzctfQa2wJMW8/
9VxjsV4D9hgTMa8CYmUV/jJRdCA2/BkqOYsShX2Tgaf3zgA4TCff10LdW28Fs9H7VKgP7TTKWgsG
a93Ufd7a0atwfs7r+tYQo6OPxOHt7iBbEBjPmwYFtBEuN1JM0Xex0QX2MtAvNud+A1I9BXQz/4bl
8iMejENHco3dst9mtmxGVvsWXZlnffSWJNb77xnHSimMvLCidUs+y0tAF6yxIfwYqq6AJGBPgox/
9XlEJeYdi0OTiIkNCtXO1VZY3FbErCL3tJ5ZyZe3MGCNjJySFWDXm4ZjFpdEFUhcR2vGKjgABPkR
VZMRQaEVyPVN0p1tlhHcJDmQB2RcQmph2BpaJQUkw69Uop/e+IG0imztB6oD+om9ze32zVaRO5+n
9e8AyH8tRzlANyNnOD1WeZ+P+TcKjRrZNzBUh0Y5TSJqpTvpvH0suV4srXF0Eqs0Sqa3TVpGiWDc
q0wVwoL40spGRxWbiTHiVHWIubyVMpounuKD2skwigsSnABt6virlfqHg73FOT2Pk2fDqj4VQ+BK
5rglrG9i1EtlJtlqM4CnkwPC1vXcWZRB0gF40n2WFPuN7LOH3XWMaS632uX7s5xrdXwbSXXb0EzW
KjO4LNF6Xb/6t/6ecWtGuM3ne5Z7oG5PA+snDMO1WkSjYdaJFPDOJnN6vo9uSbmfoVzFx53N8lWg
6IpjI0KOA73wnkZFLAgVbK/HwLqKMbBToTf44gDMLZfP9h6I9NRmXFxC2TZ8VQaaelQN4n9xrLx5
8EQNn/eTQx3CMcBjMhqv+WQGCCP8VRebmAGBwwRwWzukHMk9thpVX+mnQIDUiQhmAmywaeNKoe6d
c9fvIWNd3MtzdBircYzkElBYgy6LiveRwWFqG5WkHx/GR1GvTMPqYLILitwK/UoL3vPzxluTRwaH
1NaX+P5vPzKNPTYuMRKPQtvLAJJvWPcshyn9/4HxF99ybAqm+NkcIA6+BTM7tOXojjEZ4RID4i9Z
+i/SLWvl9IPO5tL+O6Df5OBvMNCrn4vxUq2v0p/pysd21a6UAMrWRlpYL8HjTiGG6vRsfwoh6NfA
PhbfDjJBOQZ97eupLvNyqwWs/E+gl7FP9qFYAsCABbb+MjAhymFzJRBwevB1pEbryluz6ErKR7qA
4Sxmnp9BF3NWymAC+v372MZUbUYzi4IuBrMYJPSeqZT6/1lGrHwmFhNSdHY1k+LI2feM3zpb5rGU
5urAeyeIAFsaqILAZBnGdSOX7iFhc3y+HHVG2VWl4JLjhb9K/e6AdNF245m8lfivqa81lltGDdXr
KosnZeg/rJp/ygYlBVegpCQA30suojSGuGY6EMTLabqp7zoYEzltQZhEiIUNlotpfvaIKyFNQKRr
iTnQ6HbgHlbOjfZANwdeMD+NAxY6cOWRls/yNa0eOsTMeyCRibkMrZiSSwKCdkgpqwEASbtKjugt
4K9k4crA336bjKDbkgz7HAuUdhqYrojrPJS9AzTHpMfDTcJbVU5REfQ9DrfT+G/GQneyz1hNoIYu
4W08BXLDAX07iUDkQ75yiuYMTux3bSMqee7pUoku6RFVf85/N5ZvnGJHEW8tEsuObbZF3IAfOm8c
CwdnMRGAz2PdcboY6MOi9AzMmEmZ5f+OU+evxqpEPX5KLkuMt/vEd+uYkY75VV7Sl9wlipbIeunI
l/5ZLbNtZNx1UoJUgVqnCih/QxJnxQ5rb9x9bAwc6vpfVzIwuEe8vEQvIsHizf6rIW4z7Wnz/rVr
3cUGt1YiI5j5IW3R5hciiiwCnDkPlIUiZnjI5Ntx5D3D2qee4zTReKwSymB9lzE0rowcldlVd0yL
P4ud9jrRq/S5BK9mWAcYVyG8Ig+nSfhNGv+G1ysS/y/P3qNUHQttAInMFhMMbv3/2hdSD1sOLY63
O8Aeh6SxqEhFjC7IQxiSGMUkcY1DH/zGmrAgxfmFlCq1vyzzxOZ2oRQk7XMO2jfnTmK0JcV40khd
1unB5qArAkp7v15xtDonjckbT2FQIg3Fk8+2Lu9cYtxR3KO/ORGGV4W5fqFBgoLTjAkVFbbxspXF
Lc980dFguJUD9oiemv+BHhvG19soBOTmhGbkilifua5GE6pfKfpT04QZzqTfk/uM8m+NG3u3tJoU
YSq+kvdUNkpOBObiqxdIFFfbYFY1hTbksJncg9s8WM4UFA748uaPf8156JnzFIUxkwYq5b3o7bRV
qv6wfk3KffzO01nPLc8Qd2WI5Tlu7a0XV+YKgm26cNGb9f0YHlsBhHHYp3RBh/xZeuPlzn1CYNfa
9I1QMJbb+hDo50bB/xAA5rtFShkx7RTz6E2gFgchddtllTIzUiMFBB9Rc/5lu3Z5Wa4ODirYLfab
bTjbZj/9XmECYKMRMXb3xzUdlLFFGxRhxcHoPc+ayaXv/oIUKR79M6L8UdJG0Gomz9x25faz0xa8
aVjvqQyIn0uTfTXROREhNlzGda9aeOaj3P0LM2jFWr/Mymz4ZYAYGBVDh8dyV1fQaYe7TStY+qZN
i52daIj9y5XNMQAAfNIeEKHrqyDfpfIsDvnvQf14LYblpyij4MrFyg72tEugRhBIiWfOezU4HVhV
KhPGmLv9LngKeMSI9WLlpt2Gn20NPICtuP17KVVqx6m3RGY0ug11+WoVsOxIqC9vMoE+EgJt05c8
NPGpSy2hOgPKpqWZQLWlxuI2JMRoc2SKzAquR4+SCf35NVPZ7wn4T+2c9Uhmg0RO1qT1TITfFdA1
j62qAFV/Iwqdm0pyFaAQStf7V8c3wIH+i/obnhY4HwmuVvEpFBUO3Q8OALbC9G5n1sPeEJJCon6K
T17v/+06cvadrFQEdlFf/Fwl3GInLq0ykuzaNmYx+VGwUF/aTWYt1FRQQBqF9SLYa/3fU7iYawGQ
ooJ6MHwxuwQDfLKcizNAWeSBrFUj48jvEaAoG1jBCNCC4h6h78Npr4eut8IUazPbAYM/jinKvWe1
BwXN6o/orFE5aHQkY41eDrHIqE9J+Inme7vRKs246KPHgqbjUTp7kHbEiRn+Drh2k3NJGlUQdBeV
YdjEhDa3bK35nsURxr+4ZV+4Oa4hZivWu5e2Abr1MqNniUwqR7ptzmfXDVo2Pal4MDr3okPVpzad
maXXRvgDX21KgbCSxx/dLJvema3U4VMqgi1DmWAxcwVrlr+PrJZDCHLMyWJT0XV+zB2C4PdOsQQj
aDpXleustFZPi1d4FqeR3XbU+/Bca8mUkymY1Yz+MLTZcRxKH/fx+O19y4uI8kUyDIpEAz58+4+0
gZ3//0CzEAhYrIDwQuArU92UJ2h6kTTeZkegnbF3DE2tbsKoTO0DaBHO0zhpJZfvSB3SQDK3u8hN
2G/grFguoMC9ZaWKIA88Y22u8Y5tMBgjcuSZCaHMHbp1tGokvsp1qWqNteR8kzDuSwHtOuwyk32C
6J7wIoGu3/Ia6vZULHTdHi+xe2X/hmw8GqgRau9Qm/xo7cCJONqas2GE7zBSNXjYQk6PBV3yD+2J
sM0PqQXHv8t5yVQf5uNMemtQuI2TMjCALrPVEKlYqEesWviwfVTWTO/dzY/8MDAdQiWyX8AwEJem
iXQ1PJ3Vb3jbqGgsRV4lige7nehfu+RVL9E7OtwMNEzXdlsM+TagYyG7IXj2puI9DYuo4XOVJmdd
Q61R/JtYl1+ywLzPsL9hHep+0b+sIpkVrEgX/jHDAXTtwpBpV9gNxd2jXK0MLs/2cqLiIJasVfkM
LLUlWzu/SWywi5vB3DDujpKZPgu/K82nDR1KQp+113Ab0NHLFSsth1+LQKLMMmDT2fl0KooRiO5p
ULV0FwKKrrmO1apgK5pRPH3wtfljHoM0pnHCEZpVu2juQZgwm1r77uSnEi/73oIABoFsN+RnebkW
hgo5a+CdFDkS6FF90F2wUHsvuS+7OD7zDidsQyDzR7ow7Hz2aA3PUDxw+qlbi3iJzaGJLcbpmXTO
bJ4Mf9GusOMughtqcQ29zzjazrhSgAIesGXsSYnWbLV+dq05sT8k6dO8KSc+rxzWAa+NBIOKwVVk
rRug3kVO3kb1SwVgW7mklSYq5npeqaPJALfo4D0lS5Xz3R45/vcFK6CsIqVqCfleuFfsOuTJQEGl
WrEGfBe456yGT6QLU8rbi00qO/cv1VhDCGcl1C8LZSPSLGd6NV8vETZVn6lFiVRlK1If9N+VUqxH
Ppz44dZofFZdD+ODBE9UA0fedtSUNgMANVeI4uk08e/bHdqJuMyZTQRJ/j8Ra86K2cO6kzFewl/E
z3bmd09FqUkbccTUOGMraj2DbyeX3FC54lt33gptOZG2705kqVdWdqkg69h7pX0IhiuS1gmcu+6P
hptizdCWx7dYaaaevC1DwQSoYIc60AUeufo5eH7JS7WLNMGlSoOLEao4cYh31eWy8xtz1HMB1S/Z
NwSiiOPN4R4FmTs6wsxldhjIr4EBTbzXfY6gcnLDty22QKCycQVwDAZkOPkLVXZGg8rulqqU4wAW
tKSYhd+Gh567Uvu7pxi0r5ZhfwRqWAAFmvy6Ce3ZyrU8hIFrRJDY78Gh3xCpoUOchblHZA1YWkm7
dDXcUEgNsSKkS2MIRFssOlTPwD6RkXcfJDs9M8rchSZIGwVP2MswlAMngxmoVSmPwaPPsEI+QCoR
qmQnd7Cw7Rc79FpHjZRTRJyQf/Mit97LIWk1HFSRdt7bXtpDu48VQiyHKMQZ+wWONAkf3JFuRULI
EwBJOjcXRQ0IBMZhRhojdNxfUhmAHNj913Cq6rR4wLUhHb3SEUzWxFeHtwu7oZNG88hTL3k4gUpp
/4Kob515zzsL8jIhpUvLnXJzQdbCg6sraBJlmCoa3rY4CB88aAjUsncPbpJQvmaKuGHP4RzZPCYp
MK2cPOYzQw7MrUttmCucnWqRHJOE11tTupkb0lEltUUhu7eRqTboEx/r0yy4t/xFMdOswYDs0DBB
RB4gJwuS+vUTu2oPu4Xtq2Fph2mtETOhsl56WBkFv00vDrR2rFsLWfHeeCc6gCCD3k29yGBR2eRr
uQoGh6qMbQiwqgrkFFnj8Rf0cvNgF8xhk/MLa4xlo+YLe4CiTKakeDpeER7r8v9Z1piJA1Gd1fW/
vgOWEWCFj1aFCVhg+nRcMqoebJBiAcfZN50b45Qh5YMfeeyM9u9PSs8NkPzkMzlqAW3lUbxIliUj
3vdmyNsxCBquSGH3hPAUo6U2yS0FsF4NwDDQUPijhuHed6BHAEyVoz4ZFcelGPPjhccsoc1HNbcV
Ssq4fHBS3EMtTZ712YLpGO7nlHKyTOiq5+F2Ub/AgPhmiGuYQrpjv4xRwrF5hh6fUZm6N4HTUgZL
o71p5pNsVwKJ/ypA5ydzULe9rDwJqLadtWQWkchuYllhVDkmq38L9pEQraOI+6zkQFDhNofv8ITy
1uGJBzLaM76KssG6xFpevabPffLr6aUNTbNou1R7b5xSKd6nhL5OImMcF1ZLUMKSQTLbBuS+fPoJ
E0tOTGfKrh/zsqiPBl2DP+QAnuomSKphs59IHzwJyTyObLUL0to5jbDoKYx7uDRLqdw3XHqnfp+n
hSwwtDBKAJlOKFJULXCwodtCHMWyzMJtKBNfxP7JokJoyE34FcsrzakRYXQC+pR88eXdBsX8vqWJ
7AXWnlnUnl2HJezkdjHd9VHj1kDO5VV48Ny4edIjhTFpUYzNMLtzGsuYLLh9Qc8Jji8+8+dIZNFl
GkrRj/v8+X3+D5drFfABqGy94Da4PjNlKBFjzNA4xMDE3joprzXttledYCmQQSpUTSF2inqzDuTC
i1YfALeb3aBSUCvysLQZg/1i8dWIJb/ViBSLe2DQtBXIXh4AGYrsHaMM+IvSHEr6kyCPgeiEjYZG
57jRagY+lnn0FoC8ZhAra+EEqbkAlh6GHKbjnoKTlr+YzBJTc9lJCW7DRk0Ub31aWht0i/OlYRDH
gORjceGVqQkmjZxEKJtBS42gex1XRovfJjdxNCDYVz7/+zz3HmnUHbW1yPLNuYZXh6hn4awH2gTg
zo8qUANa1/nzhAKopH6JlS066rbqP8Kdg5SHklUShrnJLJC8h30HQQdk/0l94/1k5+ti7WJSEK7c
O+F+/aMnuC7iC75R8zx/0g4VoB8+0Aim4ZKWL1g2Gl0CP7ngpwzskrZcS2v2QZnspXAzyUxTqWu4
78CdolFYqoCboU6bocjm+HeDH3LsexqXHAO1lLQWpGR2k0zTPLJ7sGwq0SDLcR8duAqOrKZpQ2Sx
OuGIxIuOThuX9gmp5zpcRrTzVWjzpT8aEkv0qdBemxwupBdJQBDfhfrmiGNzWpSR555+GAV6EbdH
RqD9NdWvXwtQWDCQIbcDaLFP8as63bPtBgMdgnaPMEPBNvEBW4IAwZxej4gTYwtFCFnH3ZG/a55I
DDCM0h5375ZwJipcNg7WL0w7i/8T/os4u7jOHbm61Ip+TbULH6mE3FZc5qYbYXx6rEjNM0z9KAXg
jrJESpAIC1u0BJ3Mx0scz1xOyMqzfrMwM98hLLvRnp/x04g3AUQPUnV/dfKXA8Gc828VpoOLay3I
AaPV7eAyODlLZGw3HXXGnlk8SdMptsHykYcCAkfxsGvYeni4uoW2kWwMUrsJQQE+Nw1Wv7HuWEcN
6r1XJ0E1XwuEKtczRK7s4bZ76rQvSHqQfkkRsBuZl3wndf6fq/keQGS9qcWrt1fKvsdmdlLZXZOL
BiNwbFOMX10SzFFePX6stXD9ll0XKYf+sC1ivJkfTN+oCLhoO9EypnoaRIoLFLes1UQ+cRCGg62U
Sz4jdJw5KjsjvJTguD+GGn9MY14KkJn+sC8IMYOfpXtXzoWdpYTpEvgZCN1CIvgoPzeB09UBjYaE
YGOkYyaZWM2uSjfNWpibLAwRNXzcP5WUCZLEatgU8ioe3MuVemlwk+w7RhtqiIasM4m9taRrkGKw
mV4S6heU/S7+RBJ69MWH8FvibBRT+7Gn6FbqYYFke30n/UfwwXme3KfSmyKyQew+4TT7mmPVerG4
HiFEWvi7dC7rwdrP/qbeXlivIEgDIvZljRpENpm9Wti/8Chnd0+GhDWY/jigx3zO6XUFclX3QJ2d
wkzaF0vKzijOM4FJRjnTLuBCwzgKEKMOvAhCn+IoveAImH2P3eg6B6jBpHfvHjga43eiSEFfdq9i
EmzpPHD6Iiq66vhbFwD7Vz8Zv/w+Eti6RJAWLtcEJ/UgsukQOa9cVYBQJrGOqdneaKyDRki0kQyX
HTscGEohTyf9pt5Q/eWI/GIebTpb+9wpvegHMRe3NU7PblAr9LLUHStbJ7kqL0dSJM3q5+tQonHb
g2e4grUmihZ6z43XGD9wKO+KorjvNw/CLiMTT91mtI6nJfKQpR0C74kbq/0z38N9bcCBUPFE93kw
xfYJM36PaNyI8WMEc3jF+fDjojJ336+eVu7+ZDMrsZfG7cd0XuZ2NL9FGW2UbZiFVvamvJHGGyeP
uC1bQoy69CfCBmWoR4M4SfITO4TllBZ4ApBzm3MOEoer8VB8xxHqEZebrSLsmyjuiKJhKJRVRCBr
UKjh0sNJePzuV1xmYjmSyr1mhAeDJ1splmAxVEVe26crDFwoNwCA5uo9lJ53c20mjn7PIcSk+eCT
PtqAdCJ85Z3dYMH23/EWZ3Q57rW2ur03Ne2FmIGzbuwR5sCMkAlMdwvESwqj9XmidPD23YqN7V2F
aaDMxD0PDQIBEpwyDJefbI0zD+HiefaN0fPrd/OuzgPisZejF4ykDp4C2+Wa4JCgwefU2kJrtW/W
mqSNhhtjsXxIh9H/W8EqF7ROhBKkzI72mD3o3M+gTWIcNDziZ/s+/IvJEOzy4X69iALWRgf0cdDX
tBg0f77FLIqyeHkFct/jJCDbMBw8inGLSUK6vTUKfT09g5c/Yk7eUQVZh5DYd7a4TnE5jadPk6EJ
Ghk/NrZ5UjVx+UI9dv46/14f7+avNLdPvX+FHk2nJrlo7Oonnb6IXRFjaJg7gfx9WTMeoZ8DmhrM
KE5Dt4VG2mT7HALoEQBRnq429YgIKb+vPZnFBO+1ld/b8tFVnNum5C2IjNdyYF0JXSneFiDBty/5
hz3XQ38k0v/M9xmu5Y5GXVy4O8mvaHrE8mkbsF6bRKCTNAD52H2382XnWAMNYi0yNub6tRtu8geM
ZnjjrhBsRcZNqAeGWqZadrhVv6f0Rtzs6T53UpDVQC6smCFRTejGXhT1Zp+Cw4S/hZEMKpxIe8NQ
J/r3RfHwCcdmYPrXG3tHD3Aiz97345XKwoEPlpgLL4ckbAQeCPJZIVrCvfPCa0Np+Qh1gcKVQwEI
O3EodrXdIIhqTOHvWTv3Vmfgtb7W1wW+161QVLSE95UWfz2b3kl8k8V//kF60vKXpsJSviaGW08a
vzBXGEjjIsO9cdxfQF3YcG0vPJ2TdWA9tUT5wB3jTtudRVZNq5kjXhHKwfJP5W4JqgRCuzMCIMuM
DiiDz/R/J4+l3++ITnSA7j/Y7PXDY7+QOYG1/9vX62JJL5K5FwSyYcqABBlhm1anBdYlFyxA1WsL
2zqJBKpeSOoASg0O1s4U6rEiphPdC4JhoEmFdiUIr755KScbBrKcft1rPxdIP4t+fwPJ0XMjJEhJ
P/O4zlMwMTCQ/JCwZznZxYK+8zhaaeUBBcZoBu7ExcQs64xw+BK8dIoNLzDxHpb3I05aXIT+thbz
6FfrXxBrxFWdoAHQffM0wzZ6aYriXi0jdwOkK0AyJJH2II4fMCMmYg/Nk/+GKtMQxde8VrosNtEf
l14MOEIC24gfxbuKwx+IQ92VlHipOVnQBrAK1qc1xzVX45w8YN3W80PT62jqDiCv7Td9BXgHvyJO
7zgsVxQ2tEmpm6s3QCikVdhpiOb3NlVU5uoNXno2eo47x8DBlwUMxJdP+nxiV7yYe4nngADHiSCX
ydRQHLuSBRu7TFBqIVcUv/54sfYSwFulQuSnrv6pDJ6vquYBQyaHyWPthpuyZytTxlLl3vZ9WSUR
PSXhvYfIQQCZv4LRvaihbLYHl8J19DRpd1Va1O479eQdP0LrUJooehmKUC37R3QkL4/iA15WzIdp
yphWTiRQ8VwAkQYe0weRIl3qUt9ttFC4gJuUPFaUrPoLr4G3rho+VbVkCWvV5afMwBIfU7SiBM0U
OZjl24Y/OpUWcEcVONK+/53rMNvz9RssSoDtw1aYXuAr/XuQB8wsxwWOPT3+OyLdYDadQLpnvGuz
G1hSvUFlntW0Iqqhk7YTu6qcJWjcfcVaIETi+M5J/zdjQekj8KkhtrGH7luKYV55fOx8yoBQvYq3
j06gfKpOYaCfzpnsF3k/fiT1/OkVZP/T4p3ufLyyvVFZyMK9yaKqj6vVUzvTQhl0MchYV2AjVKmm
ZmnGAz9FezhRvR80RMsEGOF1RbbVk3zSDf7qss/3vHsl8+1DkiYrDMMYmEhU9QAJkGjBVDXP5MmT
ZuvsKP+Krpe7DdX6VH67seJN+8/DxXDyocG/G+n/VXJFlqxfsrxxJSA1XHX7pSpmTTywDU1YqaLS
WmoQm2qPCMlONqEwKVCN5rBWRnAvZOcXnt5SuVSTfifQHE/tR9o6gXlBhAzbLaslZfTTFGWeGg8I
f+G5Z91z26elPOtytOkSjaWrEZyK7q4wSjQO8K9WP6CxFJ8zUpSO2IBTJVL8jZwfEs+/Ap29s/hl
EERLFkgl2pA6HElLeKzoSWYix8SmM2IvFzjFBPLSNtjywF4mn1FWnOKD5KcIjfYQqd1zYnkS9Ial
974bo+3ytoUUys7T06WxDcj1A9IfGSrwDdYbYhUd3R8BKonaUzWjDQG30ZOc8eWtx26R5lD2JAlq
ZzmfwrG8s4OzS2OP3wcjtv4USiL3ynk5LM/nbXmg5afjmWeNW31DBtE2z7PXT2S2EHpb6CuLwl9S
0o28GmMQ266qXvGTCQmXKXRsAu01pcTjdOvQ2b1RoBJ9C1Y8fVIU08YiCeYUSEzxGRCdSoF2+oNN
Zrd3DBYpHI0XCOCeqnTH4sJ5X6DmL75bv7TFq4kCOBKBM5k3+N/jxVkYcvPNNMXMuShr9atXF0eV
I7laqkv8eycs7fZ0Q+iA7Ssnqsvvef3eZBATe3588cFBd2lWkOQ1DfhDZKjgquI+uFXJRg5wrD83
7nEEh5PlmB/HS31+0xuhPmXcaaAqCztjhTTGtWAOrtYtUv7DRN0si38nJ2kkkPNMChDBW4hjqxIL
YhKeKqQW8STpkNkqTqjy9/Vyj2bijvnEg6QV2ZM/NfrHMFugDtCvNm17V7vnaOfIwozySxRXsq6j
X6o7sxpkmiL2j0ecpAPBooAbZtcRe9Rlz2di9gvhEjATQJ0HBiX2AqRn/Z03qkLqQliK2T7JagFB
XX9SjnLIfZmZhVDKt2L8TOo/65u9FhtMXIlqMZCdfcaR1/U8p5vU5IK7PBgS5W7u4GJsr3nXj3+c
BBM50bPXqIDb0IXfCslBsrXW978pvXvbDq5dIWHsk0EKDiGnVyPZIc46eXuHAL2lJAxk3rfLUD0D
/NZGhsU0O7C9d+7DbpvwUlC1KtRs/gWo69KhuFqKof2mS5zt09BUnCgM/+o3RMfS05LRMnS/efGB
15k258CpcAAp1NYrh9I5h0/m36H2ex5RY1mQnjbEcBlMLGl0mIu9BkErydZDROm8bZZuttujlls8
Qwaea75Ix7rfSIthkIDXaJNf3m5QKxLOvD0ACT9c/5HR0Cpcv4qDbnTIK3KFqAv/eY4ztHCa4Huy
smpLQ3/yI78Po3h4LtENSFI7SkO0s4R01pj2uh8n2JWEhSZ1CmvKkDYt41g2o3f2ZVWP9wiB+8E2
G1nvJNlnO6A7wKxAiANhstA2WN+HpwYUMFzmCD/OVK5QMHIQecWmzE/AnusiLW07aFkuncRlxgN1
iMy0q74hhKRWwZ0aEMIOXP5+zq7ivuMANAb34+QdSRWaGy5qITfTEU8ZkgDA1S4H2xxuUIipHC78
2WmeT6JGSuZ2FykEvGKSiOVh+gzoOIUClcQgCT5ALfAdg30Et9UGqNsypDKCoY23rTCBeTqiB/Bq
UkOSTjEYNOI4lLC2/JMwgPe0E9Q5TTbcCB75OUZWLgxC2/dN2eA34NbQ0QSeDcUj386PFWXkxoP4
eU+9pcgFbDjoBkcJ6GF24vqBrBPTuJ8RULS55zgdA4RvhqegUqCxbio+/JFHBpp/oR/UrE452QbO
0T8aPwr2p7dbSp2uP6THK1yWFLPMZY/BcK5oEPS5wmGKcgdgItUgY5mDuTA5vM+6rguyHnT7RibW
CUma0sXJMNb0lPoebYrcQt0fCcvZWwrWeXy1CZ70u6AW6sej+YuhGMAiXTJCAV7h+9qeYFE9R4CE
OA3tNljaEj3/wHRGeZX3jAGt/Pe/AmFFuDwCJldIJa8K6diBNgi1O3sjMMMOwVQSC3iElZJCVwlI
IHgImiwVBmNjVWZPrJN7mqLsMm0gePUqtP+cs1ByocybZZ5oyCkekBE/HY3sfGU1ZYlBZI2PwEia
43tmu7sR5b9FBIQsD1hOW5zHz9Zhx+586bgXj9KnSlfn3Ckfm88wYny2aNKz5RnVNemyVLVZ8JxR
rzMfEJOpd0rOdhiC/CiIXb5noh3Rm/rFeBS7LzJECHd719THeaYC03gfugiS3FctEqtWU8UpiOzR
WVsV9dNw2YrJgtZiLXuAFMTXwGshc7kDsTNQ6rRWIBv5JOtk6lyXQEJH557wKo1H9F2uaGwW0k/R
b0CIcDfkfUVYUfAZtaXY9onQoA9JmaDJT9gYxPLtRP+q9aStA49D4oxnYZeFa4qOHUZu4O9AIV87
d0kxWoCHsSH35e7qAU5SM5h2r12278ujIIhiLTnAxAfkrtUr+CNkhdMIlun8n4OipD8eQGT8qnO/
3ak5DYKaC8B3AWfQMq6B0TlSgoebLWlWl542PfLCdF7mEnk1lECssDusGtjRH+lkHp1Zk0oeKcQg
RBxkCS1xiBxrBNx39CxHtQi34c7ncNgOH2gcu/NqktJcfFLJjShTsy07VUjLeuehGec+vIrCoMuG
4rVS/gBLbAHlI4mMVoUYq8f5CIym+lZ4VOk6aRN3RmFjPbVmGC/n54JPkTlfWb7bh6Cj1cTkORq1
cSJ11j1kkG/c0cpEPwW6dklo8YEBH3/nuOSoBsRP4hPCJicFZhaE2+xuOdmTF8H8hW+JSwzjaJo7
5aa4V8Vdtdw9wNnntxU7fMY07SxJyMDE489TMJoXIrKWk4diFXbAhgbp17iexIuC3MpYC09TWuKG
2wt2VdBZmZoaPkjU4MakueaYtyugBniaOURvce3GDR8yCOWhxKlBnklZ2qA3ila51HyqGUNVV0aw
ZHCGj54LWINPmzi903pMR8aKkDjhoGtfMgmIk1+FTyAJw0WCpzm2uaM0rYrGDob3iUNEEUa4U0AK
vIOL8vtgXI2Fcacv+SVb6/6ycMWN4P1hoST75x65lTOysj/MqusXZv9spFjEVMSoQAY5XJywZuZM
B87rlJqkd262LEawaqPTZlUYwyp+sb8FXiz3daHb5wOWNpnDR830wBq9Bs74m4HeSdUI+Y/1JlLJ
dOAB9+CX4UyGF0Rl/P7M5VzReUqItcK6Mcwwxq95q5MFLeMNsSPuVKRDzA4FpAVEy1oVGrxV5i7r
v/cR/fIehq5d4i3T6aJm3QA43gO5eR2l46vDhvPDnxWz8Go7N2r+yMd6OfNnBd/U/8X9P6m205of
AbVn7ut0PvgX47lCtpTZpOoWH7qjnDMxfVYFbwVwjDWvA7wC1mRyRl8GhuJ+jW5HsmFe9qTypM6O
ILCz+yWwsiirt1LygDCbY/9eW2CMrln8Xr8m/wWxSTzYV5AKvFpTyyBLEWpg2mNJfnPfqKteuAHi
4KRbHwklnPocaR0dBppn1pUTpTDxgvGvqqTHnUDnxRjuol9VnyjoIRcjT2KZ3J4Kxmtaf/rLMleM
I3cO7alQa4zCQRDaXSDPv0mxMhkrOif09KEDH0NGwpRB6AIeMpNMBlBf7atmlm3BoSwP6KhNhWiP
0yjSGhPA4sycHQNQy21yeuh/mzGv7+Rc5BKsssvB12kb64K/UmZ6/bFAz4Q6HIgWBXc2xATRxbhf
76EvuHMHVNtP4jJtQjNVhDa1XnEkvfitet5BW70n6u+t+OSXTA34J9w8SIvDn2Cac9ClMQrQ2mzE
e9tKUFs4JWCfbKbJr2Ecx1YEenHB4xqEAY+y6wvao+5dO8qncbz9IujGBE+Dzwq3Mo4SnJ9u+h7V
9rIqAwqbedSXX4aYnLsl9fUolHfhHp7VxHn7G8AdbeKPz3QWsYrL5a/W1FTczaiEEqdR4EhujnD0
+vQGBTFi3YpjbE2i7NbCMEifQew1ebdgDLZRRVOmSGLSjFQivkSfsBh04qPKIOW77YtuiF/NgUAr
o0CncKsoymyJZZIKoS2d1T0LmXluuawTqME4wSVl0exoHdGMPFv4SA3oOB2m3McFd8fBxG3ukrJO
UHmzab4QcP8QV+Nv4FrSvDf1R9fu+cKodNDtQaiz7HScsrKnV35VQZjCnRe1HdYSNWrT+gx5cqZZ
BzI81MP1DllXSN9kcx8wjQkztgQhSnTpPIDx97uKR2EQLRm1kJfFMS/8Uo7m7qGaOjhZOZ9/7QEN
AA1U+lgTKpyaGei5BP0hYq8mazyjjWEpTcvLEhdtXfm1WktevwqGzx1PGtEBw/Bph5oZhJrx+f+9
+J7xpKCwIyBZ4RkocHpDaGMq/5fl84QGlLwu0IWdOqvLMFjI4+826DH/gcztEbidAaBqWDNl1EmN
qGTxTzyX+OMYTBzmMsdkUSCyT2YIEqPt0tsqCJeQHv4Q7TXkn9nMwu9SI128hgc8jZVsr0F+6nxE
r8UyGiEM0+b7YIea1GAQIdRekdugS+TDrts5acNJ90e05yvvXEN5HCwDPixiDXCzR0WdstcNBIkt
+7I87sscY1oYK01iDK52ngbXrF2nHtLO9QJDj9peuPTfI3hzapMTsipybLROZOwM3U25RH5IpNsl
MbV/G7EgeQ1eFgJCQZWDeifr/dwUAtMcPvlmAn4esf2S3HRxo+R+YKAIoYCy9t8eXo6variaqNlX
6NuidID4ausnDjJBA2ypLkCxl+qX7PB/A19ykoBZk9CmhRqFC4+OHr/j+BU8IAa9pElcdEejjg+I
YELukXZEGSnoLX9Vygeec+a0MpifwiVHUaTovrp7FohJ6ZddMGJZ7K0lnsIu+HgGDlRBhj6WCVne
fYHRC5wpQEbYcLHY8D4zw4IhH5UXIaruVWQ1W5R3rhhiIwqa58/EaaCBHPrh6QADhNLWv0sKCF7T
w8MAvlsWs7zwXgIvFKG4SkrOOEmXnUJe5UqvWIw1HSjtna33lyV6ADyWJuickCFmJ9ZhBmL/upq1
0TxmUW7BL/V4HhxvD61zmy/TLHFVua9eWJlFtQ0ihaOqb+TRBhmtoXmdWCgJv/XP7tU/YdyxziDE
9qDcOJAAYs6EM9M5Z9zz81bcBSY87LD35JqNNOkPe7HDRcad5Hv98KTyPpm2I44ZaYXbLMbulbWm
RZnN5wCPL9J3D2u7gITR+PuPpa92/SXE6MueUrE7IzXjLpXQ0ZC17jAeRn2pkpzR0MbZ+D6dZWTr
NEtULFgbmcHe91TKWvix8qZVVuL9ss/cF3zqc1TV62VP6lUxY+AFDQ+nqd3l4GVe+Vb7mqR8t32N
Q9v0yYb3x+nI9bZLLWSbkOnqDFmlq2cv4KCQVF5uwqDvXTvr+KTYqt5KobOfAydRTONQkusdEw+I
Ei99HtuUZ5FSXCXo1fBMlI1RtyQLiQa+AbkrZmuey8npXog8dE+nvTMrHQLEw9tpHhvkbNONvi84
sNc8+DdiGd0879IW7K+RL+r5MeMOg4jSL5rcmxg9At6V0wGirRoNs+/20+/QC/z5CrfHlPHNZQGy
omJiOrooWX8uNCX93ODakiO0qBsHTxALWlRIF1Sk/96IxO1doJ2bDPEGXfuv24cRdetdZzBsy3jn
VqVAQ1JbGepqtb45IzeqSp74Cs1HwatqJQmEkT3rdrYxrhnSGD+iVzVmvGAS3M/9WIDA03Ra3cHd
V9613fOTx+YMgI0GN7bmQkdYmjGKgYVZY5v4K02uf+SzVDT1KUNG2EHpRZOa7kBWzeGdAAaVLUbg
nhgtKoalneVUNaMu49LecbyMRcZRwDHMcOYFN6cSWD9HcNmVbt+fW4pHZM6jOYXY1chtJyqxa6Hl
YOO4rqbQU3IuxBYwzzXrbvPOasJlWVgLUcm0w3SaE91z3kz6FwiP1HQeG/grend7+UPz97W7Ivze
NC91eBMLvKfr+V+/6na3g1ALevO17yg4AgysUc+dX8PH5XjxyqgXdGAaZWJDRD0h63g5LvGu4U2W
wO6mNh3IUQMNbnOB/L0gcMj0i+qXKrjzdfabF1zwxw8L+7KAyHfrFP0kOSi+/Kgup83c2Cs2AHuf
Ck2SCWCGLpdk0tFAPw0e8p29bzOwIP5rtbPvaOIJLXclFiEzrmobYBvKMQ+0yVPQKa53wW6rLXWD
cyUem1J28sJf/yybJGoTxKY4skP4ZEjWe3nts11AuEtr8hw+XEB323oZIBDsVmR4WpOgx46D5xmN
hJUROJOS4cl4myU7jZ3S7WGKszJgEJpFmVJ8sa7lBZsR2cLoUdWa85kV7itdQMvwqMRDMyLgNyuF
B09aVrvgzIfe1zaq4NcUv2hto08sHanVgnQIs0hzVRZ1PRn2AklaqQEgWzXSYHGTq7oqJsBTzTCL
BJP9sOVzxuA3QKII0KBf5OdahpRa03BJaw6V9BeghEInVGbkLLNVSeL44krFBjrDj0YHi6W3ukCv
XmG7yR6ohGEWk9CCE7HXWHpbW5qbZLD41TpvcGU1HZISfXoy42TkYwE6Y2XKeY/3qJcsrZf//ksS
MQDTA00PloNGRM+JBkiOclA0998vNpnEyPSNaJSAc/khUWX2qXnu2nFN/2IUU5Bd0zQBYyX3pPKT
YxKRVNAPRRzoRbHWC4XexY2ZshIQaMsmJt4W4J+Q5zE1Q1Ym3B7TwTSqg0Ip/kvg49OaHT5XqoX/
/OVeWnxa32BxpsKKYtKGK6SvzZ7sfGPlf9+cTM7FT5o0NxFbdfWZzzHXWjAXhoULED/5NYOrflgk
KLVY4ZyCXYc42F+kX+MwJwraNFLovtGg+TnNEqLydZ0Y4fMsa3dGkN5X/07zY11G2rmCzoRD0+RH
VJS1/hJ/YhKR3Ah7KEg/VhCbgAJqR416KhGEiWG2+p6ywBhvdxrgqSpA/oySD+XjDmpnTYb7a6RT
CDUvkDSEr7J1pwFPDXyfWTq0WK0h8aq1+zmZolb1wmXaD1WlOKp2Ay+zOfqBuUNFVvocWWwmSfqT
WQWejQpLSfuDAUeAKcZcv0WAqnYvHVWWIp+xWfpdDRe034jJ75TcDeo0G/4Whq2yx4XZdcs8ZFr1
oVpIXwjYqasIOrOfAkAGvzBLsnrN42TYPuzdtFO7++77Q25lldzm9Ny7TelTk42jYXCutc7m5CgW
yEGRelSQMqOGbKk+r16c+m0lP5oaFWkJtv+ryH+RhdW4xsJEwp81H6cSILye+y4o1AAVh1crdbkI
LgjZcjY0rhHgvqT6pV1aZstOvDuAN8Ej1BuPQ0wGxZG7WM6TDhTjdhAjYdNTIBOdqovO5jzK4Z2A
+OHlLxEqPuQzxFEyLUxeFUdyFTrXP+toMnYkh3DcLnBvbbzwMMVivpKhJ1MVP3WxWx6hbo6FHKny
ZD6Yay4ty4uMzNenkF6of6Uf2KLGTnqkKda1EmpUTaNkPcxhBQ2yv2o7zCr2tiQSQV+XUY9iJS9B
ufchHAG3CmIL+Abkwju8bvylVUx2sSezoNnu3TlTi4b+0PEq0LN1BCIm6YrQ0YcBcu+qp+nceZcI
uEFCUTxDvc+dM5gwxQgs0UH9SKr1YURGC2/+8IyqIbmxm/C2/PWokLcz1D3vpsQIdrpA8mlYxpOy
uJNPiNVBpg9gYD/H8uqYIbchT+Yrz+sUu29dNoCmfhStH2GDGW4oZ4cbcvipduDCrzDX6MH3Ak0o
ShozerxlLjffqhMH+ie7FqoS4/n8M9oq5ujUGoiuh9gsbR2Gnnax9R3m+wLomAoqm99HzYiHeLzH
rPXKVHGXaQlSezQ3WphrJT8BLNrtvaRsXfc0Jo/CoJwMmcimXxv0Q2IB3x4GoSEcBHn/M0hWAKFY
XE8zeFRTVG8ubZMWwjq/3Uu1c9khRtHW15m1VxNYDrDijzwiJCkZTj7IeYCExxdNG7LBG80+KXsg
qckL5CrK1QYdW9OK55pyTw06zASlOiWnj4d45NRO5CXgDIjlBHf4j5+pkssfSHytUc/m2u4mSbR9
1yPSnZx2m+80API4VybTIkOWrqnvED48g3zRfAgXGkg4eWk36FyXgCZ92vRFi0ArB87LxuUWlrFo
f9J6TQASbCKQZVuF9yLVeYmACSSjFNhgcyIe3thvvWkLYf/1HDoE7812QTg0Dah1LQ5HzGkN97/i
np3lkkXsrS8X7cqAMp8jMf1cH1BXhYH4qHro2lhdctb1bs0/plirO/B7E2lDAZfUMjx/VwALaB3F
9onf1Rewxy2TfkfFZt/YafWr8wTmvS/RLbDODF1GR0rRVf1PWA3TL4BgU9zNwDWeJUBcWAcP8h74
Z/M1SKjHO2kq4h1B0KhcqZUDum9HVx8LUJ8qZlbSS6xWbxgPEmHlP0iTGT9LtM8+GGTrCDevVOjt
J+vtbAZR+4vg3kW2+eq9LIMVOQvkCE4EyLejQTKjsgfpWKnKfPuWNAcd3IpvKBS3dx4r+TSx8Kc7
lxXABGcz1SsVYt2uq7DNHZu9j7OBjRlhboahXz4DTGMhNneZj8HRfgnuScVRlZutQ/U3nm4dY1vA
g9tOB8NM1+mBzwpStP3Gw2yVLhqZe6SYOraTzMEgh0mPnTnRuOrTbNnl46CKGpqjxnE/ja/58K1R
43OxNl8IvWD9xeBjKIuEXiVICqNeRxkOPa4MXKBiimISxskGyZmfovrniGGOukMCcTDaO8h+7FiD
mXhie0Dgx7KU5pJapBc1kqUd+gP6mNrYWSeJXBWDx3Y46/Ri2g/NaHtPc+3p4kecMBitBa9BbegF
BglXKTpk14rxkbgE0MpUvJRbjq4PGOxz9kjEfEFWx/dkF3Q0+siTEq9DU4t9LYSdukpRldVGYfXG
BgetkPHCRcjvMt6421l28orwcjL3k837L8whvBi+1+xI9lyATEdUL07n+zcjXWeVtPtymAyMyGQh
0I+bE8ca9kTeqGwWsL2dVAS08Gzdr1mi68EFtXwWYklNdlMlQDeKyGkGTdE8TBIW1vNZPGwtysnW
+PZlDYuQxXNDpQgNCNIMIGOqiFaIw7dnx43mfFfcMTHgDb0HP8NImB7lTxjbgDRNEqfJQMRBH1n2
xLFbelQ+2aoBk/HAhyQv74M8P66DTW+JgO+6qFKZy0OWkiUvfZRy/e/uiZrq6nf9+gXdo5LeyjPD
o2tCLZ8I3j5r7BFy7Z2HYO1GJDyDT6joiQLuJ3A1HD2VVlaX3DXiwV2vQl0Ucvu+soHiTuino0mU
TnLBja6V1T6cfZY7gag+33lnryqlMknSP7yMOxO2fGjhgBxLyqVe9K4ZDyP+SVjFfodoPeFKkXl9
UL6eLRw92OgwT5X+Qj5In1itPmVajHJfKxpyYi31AonTxSJyDVpxRJtn/Q1lZrQCKILqgrMlnTyF
yabxI7n+YDmkcnspzN48EmbnaArH8cID8pEbV7uGam7uCoa1xTUcuXuhnMlyYrm/N1Rb4ojB0foy
so9xaWAf9mCtBF4vWkx7PZbCG/U430GnraUIVa2+dmxvjXCluAInRpEU8M+OZ3/E7IjG+L4s3msu
1Qv4w4PL70Q+V7dwvxqKKudVvyg3WK31klutYpxA+Ajn0UOfHpQoyR81alAKD0fiblFPrC7/JA0M
3RostYVnI8XyJQd9pf0pEXbm59/bj2AttpHuX4lJmjwpapxxzYBkN+2e/YxeuEh3BMPlRoEnunAb
FzppOAsuF0LGzYydDPEoROMU2S41Xfu2KDMa4M0Tdu9YyE4N5PNXI/mlQeP8ZYgS14ijxG8a3dEc
Vy36n5iCBW+h93oKu4l38Z1cIo228dDYk7LMT1/6xm/OmdXXAokhfSuFF6AP7MrKKUBi7FusZ8rq
UNMyFE3alpQYF1Mo6VI1bKXlhOi1kn5OGkL23RK/pAh6m+tSGLYuewRsBAblKSnvP6fLmcCVlaxv
TN+7UJQt+kNAnx34kV8xP7B4iVIlxhQtyZnQT+4ArWbi1WkToS6c/HNsRRqmVsK0m1/7oqdyS41F
tp2OnLe8P5rxTqZKQwhvXfjQWqz3kE8DBoz4eQv2RkF+S0htQOzl2OOFDFWuFjvTSAfdLhh7/YNz
SiVIZSwnoQQMHuajAtJmc5BohxfkjUsDsVjaZb3n+Un6gHQIcWxYIrrOl0mhxqZ2Uqtn1u7ynH39
ompth0rnNq6lti1Rht7MTfBF1mKHTaaTWMmMq+JhdQkzXxUrOV7Zlzf7nW0gK6fAZjWa8wO4417+
KKnMSVj6hBpvZSPWMc0LZClv7/5TtPnVbr7hpJPm0O/CgTbTK4Ij4+4V+hTuyUOwnjgPdPHr+v5Y
5Emj9zjrLcJYhpBCXay4wvWrmLYperec8BpE4Ct+Xh5UY9lpsoWOb2GeKONjRcPD5ay7nBs2oo/K
jjfS7IkX0AP3DYKxPQLBWBm5j7FT+LxUVOdggOyausFrbSTtTZzdr8A76hFxPFKNIxM7h/v2169F
E/qvUzRpOpFX3FiYO+asHtQtB0hFn5tPQubnsR0ZO2gySl0QaN7osRsgLiUnSry4gHVKUJrz5eyp
0ZprrTaVRxRvdJsUi/8FPHkc5gvjg5KLheUkw6vpKLBnEPtrJug7CZOvQQfCNhxzL8d970CrCxFB
17jcM7K8XoDTfmM4b+pCtwBGbtb7T5ejsnIZgMtXFiXK4/q5Q1iHez3uIDmFogrSSvLJE/RsggMq
NSBIv+7rzxsHJcU5O9ugv+3jY6pfjR7zjQubQ00dSiR6VxrcnQZTG6LlTsRnoQvOoNfPj8c648YT
bVlgfTIPsmoZOGZMrFctXn5qQQEKYnDEB8MHm/1lhCOXiwktmLyVfn5DQEHagDJzEFEIBTzNi6+x
mg+2c1g1vyljVJvnYxMPIBhvDti6y5TAZ/OB5uAdyDxvKtVdiY7bWTSeRAhN/xvyexmyfZHGlVAZ
4LbPLvtNaTkbnrbVh8keCYeermdH7E74GL2E52Th5QhYauTVcHkcsg3NLRAOJUnF9T78zMYYW9fK
7Ivf8P3lVZtvIt81KjaSsGJnMue/PPEt99NLgGDbc/ejWt/4eto1YgYYOFwSVxR8oXiS/WPZ9o+p
G6JMtEQwZdW6VrdZsW3WtBdaqCEqtUPWy/g3iHVMJJw1MOL1y1fOrs9MMff5NGUa+Dck65lbi3PK
7DO2I+TgihW9/2cAVx3JjGK0hlxX4v+0uCaiizezrnt1xXjPqFUFzc5VmwUyUJEVRCSu3cS5X/7M
TczuB4h5LGX6sxqBTIz7Sg1B/W7fMOrlvlQZ9G7SAH8VB/ZW92k31f+FJypNVw8tw9yvia4Qdsmj
bcH3dO65BjDoAETIl942Wc+hf8Boi+6x6noC1k9mteIhulkpqr9OwA9SDnxCI5CrFZsrB/8aYJ65
C8uqp86DBnzYBebL65JiiFnWHUxavsmbGfaGJoSA8f3WvQxQEo5L7qW725076Bt+pCY+fKgb2RjS
SHxFRIn7lHdo2QNROVJY86+r3VecD4My3e34AG5rn+RazZxeEV8pK5TYYrtEZkxObOc7fBV4CfNH
tLmfdY4+BzPqfRlN1HVUKkQjJYmUNDT2RKMjJoBvV579Y6Yd8jYXSiH5fmnlUA2CTcGX/5xx/mZz
FTKbEu5RTXf9isoSP8IiqPloT/XQqMAK5LoKy37HssBUBjUJPvj1dHtqQk/4dVkJNEiQGwnlkbVv
40QWY+z6TxfhH/y6kqgnJ4kzuhdfuZ1O3SNSBsP71CYeVBZW0vJL58Bf0pC/V7F433R2znDH+Drt
zYRrY/Sp0rQtQqUcuQhSLzwF8mOG4tBoPtxYzJqNxjQB2La+Vwi47nHP348azdXgaCdDfQ5Nk5KG
Oqq4yxx/an86E6AduEKcpt7tNFLz3ZftGjx08O8Q1pwSeqYDEEQQMxK3ryYc80nzX3tOUNncYViN
AdKHpB/UHBFOelfEU/BbSgT/khEZ2siZs6hiUZMP43AJeeGUZRpqdtzEmfEqXwju9ITWdTY3vWUM
WpEPa8MR/nmiQzMn6/doDWayFppa1/nrizmjV/rPSJ+N4DfjWNDeNTxQNsX22DoISWn/eCnQtBw6
3SWP2M7EQqehwcMUEjsH0dlYR+uHGRDd20hJOGjVibISuxg+FwG1Z3PdzBZA8oIJIp/+iudzj1vF
Wttj739COX8n0oG0OnwxdBkkllH/vaj9afQcSY+U91EBzg1lnY7dI/UQIrPPw/xMfN1IfOM/61na
w42ae1yZYr6+gjwoYz4DNFhkK0KRMe0ZRjCk82dybu03vmZHU4eHuYWDj/MHTWWMw+LuDS83GBw+
/J1NSyTGcOWx82G9YCtUGElm+QMMPGEv5xrbqQpXTzx4TZX6BoPMpniTg73M8NnwOFptzpN3BtN0
bOn2FaJiMwFK+isqOrNmlyBDP28FWjJpN5kHI00fNFkLVuBaghDhrdk44iLKTrTKn8I7ynZG5L+G
3KezAIm31KHxNMVtcqf6yt3wRFyppJpmF/g0EAIDhxyffoHAfb5xcwEwUEbylRg6rgL+/vJhF/vW
IeXQjJZYn9n6E0HF6FKBzQOne68cCM3GKk5m+Zuksiiy/FmZOYwtNn/xkYCM9LtLDkBOVD+p1Ihs
UmsENGyzIHtYvjldxJdMUy0ngBgT53nIWcxY+W6kBKl36Tflk4nyD1QahPd7m+Un+/VcesSgPztj
l917EPlaZJEwtKUNIh1qdNq1zuEYeeNIL/1w1kkVWadIqQeXl3tJcOnMRIvoKly7v6GwwXtrKyXA
vag3DAUpe/V4rLGij+ciQjSEzWXecTBo1Phf+FG+G006AsCA5HdJ+wUK99w/SRqMdpSRZsMDGGFi
KJGADJqfwkUC1fLHJ5/EllVnv+MU+gjROFKcmVgolHs8xB/tlm9AKBgAipTUx9xkjEgNrIXsxUNH
6MQ3H4BF2lievrRWBvNk6Vs7oKibPp3gpf6BWKXx1yVK9Aqkcrs2t3wHnMQqjIvGfUfCoKjiZZnS
0/L4Oh9irapoZM5qycsiIbuFbp0fIF4BHY1S8PjN2NDQoe0z27fsBfCZSHyXTP3P40X3rr6u4lmi
2SG6lF0qaviI35QheP6mCGf8ynPTl0zZ+cSuxl0u8R45YZo+BZPVZyE59LFCkeaKJUvK7S7C7slc
auABej3xMf+ibbh28ehgQ1V9AVo3zw+dhRQ+6YbuirOROFpqwroUaiQ1TJkVyYB3nST1KNaAGDU/
qDgpU8cfMlFJnmRyLJ9oRejXVTZ8Nqdk3zb2zypy8DDlwvvEdeXNmda9CaIGG2wwTmDIzKKlYcvw
ABCbGTeXN9VNdrhz4jaF8zHornzH1WWLpANdhCQSWDJjVhng3Mr9yNmwFW3GNEelz2vR5JhPppqA
YkZU/GaLs3/eCQ9SKMu01vzNzOpMylDASV83NXaLmYIxbvRNCo9e6+68NyyreygVtJ3DKkru0AYC
R8UEv2zjOG+bodL5kzKOviivxpQ9SWWLyMbphVyFaIM5EvA2bGHD+GIbQfj0G3VbTCWJjlbYeeVw
ZvLX2CTglIk1RX/b9SnF6a6p8eQXm9p+vZ1uF0zK6XPXhx3QdF+aIyBrp2rcaHtIyaQmQFd9dDg5
D0uXLnjxJA9U6LPZtqcGDDk8+ki9hxFDNMs32tvbMAF4sMT1Oe5T5C6UTLGUcLQ2gvXr/Ho8O4d/
RlEX5Ow3Of+toQZKKDfxgnX5H3D/6IAw4woNLaibbf5478B/gQPXZRdL8A0e1FtKsfyHNSF0g3l7
xP1yW/nrqXSEMvVWkXv4CWVof52Nxs5tsLLTxSCQm1dLDORIvTyDvrDS0mPos2WOfIf35kALlrGB
WtVnWJC1c9CZvhOYK1wlG/+EHMU5QdEeM7CCjw8HwpZdGNHp8DlYzwkn6MjaY/5+A80KvGcG4IZE
KVCm5iZYCbI+Y87agx71sWmopa1ZYT6n6VKyrK1XeF6Ml9fk4tyV3QOlXDHpplgTrl0A2cxE5kHS
WDOPqM8JBTjoP4k+SsPU0m78aAtL46vrrISGXV7LAltlR0fxwjry79Tx3c+oGb/rhETfwWWBILT0
Dv2y+Tyk6lqiAhYJMuGwFkINlcwyvjldH2PnvQVtkgN9ibNCWPK73pLxuq7hcF7LEVpHHMTXmyhS
UBwyBxpNC7voa3IhJbzQnjhauJifnC2aYkq4hN4KaicSapfbXkacU6AdtnwzbKQor6H368+NBFNw
a8JfTi1Jik68NsArbRLzOrN/TeLUzqba1H3uJdD6PhPpRbYtRBm8RvaIl0pk3wg57bEsMzsw/CbC
FJBVOsMga6/J5fl2PGK3KZ3Fpi3iU9dZfu9dz6mf+XGf77E4LUawV4CaamQtT5iNzwad2P9BEqxE
r/7UE2i7psNdZoZ+tNbzu74i9mxvfGNSA4yVc/mEKVY2N0ncWzf0p38TzNPaSAq8udf7VTkzz1ix
NzngDK5WSyMyvlZXxV+keehrbCtDMkCPF013r2dfoGNdvQ8Q8bNXNyIGTHvZEHJCTjVLutTMO4W2
ACMgsaBsI+3dcpI/6cC571UC7iLwGNuOa3ip+zTt/cC8pvgVCJsMNHoVpQNF7yBGrXAu5LuZXZg0
NUAIkkQzbkNJsKV1LeHRZ4Ffrh/9lZWm4ZKWqTQEgCAe3thYGQiXOrAhhW7Q+L8HsTcs6DiLknCT
aSO3Pl2CuBQnmEdZh+NVr5sCmyU7/p8c18e5KuokRhw8IRguBfsqfiaeaer28ojWz7GhLP+HJKSJ
xK17cjFT9uU3sowyhHqGST4DNbFKqGVaiI+xVD/Mo6rqQdEOXkduFDSy9t+0ZOC5Y4vRl1vil3w+
LqqRB1609n/RaKl4yB9jvl874VgMbg3iq8Qj8e/PYB4l3oIYjRpu7ygJW1oaUQQhrPYxIiLgIUmy
VjQiApZ67Uf7P/hizsLVDOG7eFHAmw00kBIEf5k1mnAeM1Idk14Afuy/EAfa9zIJeK4j9NGV+gTs
Hb7r5/KCCI0mauklbzGlchA/er69dk82yFsByWutO5gJsMKdNx6Ml2xRNx1q1y8AKCgFBaMe8w3z
aqN/T2/Q6f4nHB5WG3EiMMEPmu5Ll3L1N4uAV88D/GUDgewSBkKJqqaWXwLgy2XjJblAofKnF73o
QtsQaNkovZSuKrv+IY5oT0hG4rT9XsH2aeGJwKZUUwM6CnWfQSONs4S/GCK79rob9g0oqF7u3yIB
T4vinA9CYlZUaFVoLaOkVM7fgh2ursZg4qBAyw/sYeMEhzRTdf9VQdkr2HLwh92ujoTjY07gNn65
osacpdMIedjBj++wThMX8nhOTOUmMSAMHi1JuClUf+gQGXLyzoF/as+c3VdKPeEk29aRSaQqxlWh
MTib299v+hOoEClU8kk4w6B8eRZlFPiWPLpbAMur60SdWjcep6pXR0YmEwPBbpkKGAQZVvCFRuCT
hiK+9rVxuhANugxwiPsNYotm2NUqNdU6Fs/p3192UZwhwNi4RQ07NHnQRfrqsKh0yOahU7+sTWjY
xgaUF6GqkX8uXovl6snFEUV3JEeR23J0vglRAh4xoKT89ZJDz9w86GHtX6sFkZluJ/IsrRF+69vm
8iBIBxlB1U+Y0UyLHXx74dbPuUA+wWx2xhexbdix5O20OnkHOgs2hLEoyFP2qUTPCcSqHZLRulP8
JfNdRv6MpzTw1PWNACnW8vYJL7K5KQNNjp5pTEmdLzbdCMkbJKG/ih4H4cc+5+HCTKU0gja820Oh
gN19zVZmVBKaChQ1mIk7dR/uT2wVRmJ1IbW33u8o46n6iZPVrMsIg7htlpIEPfkEyGOKDqac5ht/
ucQNF7Z9TYVLHxLA5ckh9C5jHCU46EOQo5EdbTMGCZRgL3LGHKC8y0jWonurn/3Fk0zPi8re6QO0
Enlxj5GUsL+eo4g9I3asNiYpM7nBu2PiraPitCZ9b3B5VSaNQ221V9Yc9WV1oGV6PYDwXQXJK27K
EFUnRwcU758yV2DzcDEgJXeVicvZM8Eryyve5TtmTkY6mdhmrtPW90Mjxuv5OztQPuSeIYf896H2
Evl9W//ckQ07+OGkV1S/HsR7LWofgxtVfcpid+XH996QPIioro/01Qhy+BxGGPN6xlqZFtB2jYbg
pIu28gAyIkETKA/DXsubno4F6lb9i3A60d5DPxiy06Ctt45PWFXMeq87FiKfeBjphZcKFwzLBBSg
9QrJviX36FMVit9OJi5aoJqEIb+NOgfnvR74ETTfl1+yDtT1tMsY2Ag3dFLNOJowiKZWylOCx8UA
kq3enZ3YO9YUQFOPqz5S3DKrfjasm7a5K4h/qpXWhdXNL0hFAFmXuCtk2mHoGlCjbqovg7UYPcQN
9moIF/TFO/2Ps4snGsp3eBdrYTyZ6XZC6LoXPd/qWnjkONfPmdJxFZKjSZMhjFJMSS3KVlUhUfY3
P0WTVaURqbLYGJO0Mur7fDjKDXoyTuDLTZvQq5VjrOM7cERzIbk610/sIgnSEJ26F4W3CtGCTJ6l
mOEMMkfYXfcYZV22kZRrYKk2hJWx9n+Es7EObZZksWZg3k/t93iXgDa6iQ9YjGne/g+bhMsLsXqW
PCyvLYDiflCk6M4LrikZZDbWV2EdTGlRvzCTOv9BEfB5MZcR+cIeXf5DUqms81QrXpKx+VBbXY4j
NRUFYaU7q/y8p+daBoLiKs3KJVPC/i/TQP6kRbl+k3jLtBCmwGsX/yWr0Z8lglT8sOqJ4Q2oTIVZ
uv/qWGhfbMJZsMRadkDzLF+H2zOmZscnClTwFDQFhB1tMfBWKIOw7miYM0QYg2+wDukVRkpJNTWQ
R8bRbgog4d4RR1yrWQUMuthBtBmAhVnvZm4WNDnV5o1W9wL0yb0ycnnHegXbnt4KZknH/oQJD/39
1spoZvN/3c5fNfmtqXcwFXKOaJmjmYmd2DKf6oXK+wx1Ft8gV0mf5W5FFoNZugf7i6uRy+pE31ZU
G53iEAKrmhiYmU1bHtVZ3F/PMV9isUvBxMy5TzkjUK/BxsyyfWQeJiILIyQD9aREMY5Aq+BRPnDE
KA5w6XjgHM7oJgkGqEo69zjv/+fcxTKSvtvSM0WiBDi/WeXp94uL2QSwjILdJqkGGcm/i2QGV8+D
ASf4EWRd6Pkdtguheoquci30xEPZnLKQIUzL05E3fhQ2FMayoYA7Tink7/j+n235rrOToOnO6DPz
JM8h4io2HqBvxBj/v1t+7QOjup8ddpHc08K1e6j0dBoHNA20UnzMoOvlGxefRkDCnQJEbCCcGVnA
06QgJGE4GbVvppSZz4w4foj8p4SmRSS85SO9KI78pGHhhwwoG7xokyCigNkWE2HLDbomm7F7gutc
d2e7wwaeF55KgXm8tx6/h6tQ8DI06CdBCE6VLVtKtLPi5ObNYtnZTmacaaQGpJmhOInT1PkYuiTr
HKfYrOnlpY+nhEZNAbNWLqP8nsrJc5QKutrCVF5dD3v9lA1nl+8Y1bDDwuiDDegijq/scMGiuaM/
HfRRzzRAmNzHgqDe9SeOcS4KgBhTATbuwNmTEvVfnYbPzu6DGcxDTXTc8KvBaI8UKixL0g6IG7FZ
p/es9ZDL+HiDmU4m9pGNI4/XJBFgE364MfnEJEUwZeN75K5l2O3J9hJP08m9lcqCgVPj9jNHSXu+
uhCM0eiaTCpwTM3yMGWmCP7LXxRh47/hGLKlybZbDNyrIOZCu1xRoiEBunQI2Tyqztkm7nxrpm0V
BlAVpZlsOSu2tUVRhpjyCIy1c0ovrL9uCuZXlzE8s4PhwzCxKA83bSGC6mm4sjBsiusCE3PMo/zl
7mx/2efrzgSuXQ95Rbuv4exjnr4IiqhoDuiMkXXURjAy/R/NUqWk57Gmt5DUiSxKdbgp1Sc8uPkY
x0j358kNRQOx8dLixU5HSogtZFRurCX37OwoQj6pCCyNWvh0myn7bfsQe1dIdxlL3goooX99GSCn
Uo6C7gYS9udXM5G9BwzoWngAlKJ0v3gA8YRRlywhTSNeryX+5jhrjpLrO0yT6F5byPOjHIhEueUq
NIx7cK/nE0Yv2cmOHqlFKEvi/8wMy9SvQlBor7BHX3zSq7WKVmhInmnQawSHUW0O7bvZmA/hTs9H
nMxfdiDMEVdN1ifLJNef3n89hp1Bs7j20kMSfAEm6hqSxv2spC0xan0iKeZMHjvx8Pj18JaTSSlX
XX7nVVGSzvuzyXGnKAPY/MQ3SoaBz+h8Brc+k7tQOk80xToeOybCJUaPe31mHIaytBB4zjREFiAC
99+G6Kgm7tLkcQ8Z8atCGAazF/wbZeB/pgsipwwloOU1sVzI8c5NGOtnGFcdB1KPfHdI20v9Olrm
uObwsJ0DGWGFxDXMjri0nHwh3kZkV49EABjN46PCzxptzwCeW4M7W52f/N/p3L237UiURzHQLcRF
oSL5dX2EH2RGP0rwGNaaLDUuBoSgqglR3SPBU8fi4vUk3vbxFpmDrI+MvEp2+5pXdnjl+TmWhLrz
2MhhOJA+tyXRzJ4zBgDXzaEjCkVsFSRh6uK+UbEF15SUsKJzo4xME1763IODkMyEWZzwzGTQ/gXH
bknvEo4C4wLBRDiyth6uCgQ4m2BcnWflFSeSjVHwVzF85RsOVjjcTtI8Pu4zWRddVqNYOEM48l0A
N2ViGMsFPImyjSTwS56GkKfQdYotQ418qvDrapCpPoXBbAmOnB9qphYdgj2e3Xj728bXCPSTDYin
eM8O8jm7IOSOHj0MG4zZrWqHcUMbimKcpXjDjw8qtZFRPUR5SSd5Ob+zaJ9x1XQ3dLcDbIK9Qy8E
d1SmKD6DMyA5joR1hrwnEJBgsqXUqYURsE3eDiRa3PbNS7EOB3IcuPLQk3G4hdeExqUMb5aQe26P
JU2VsgY6v8p8ydOzQsQtU3KH9cSp2kpUdbloiNU9IduDSq9A7MBLUE7v6ytpphdG6slU03DVTZzh
CaQLo5ap2MMwVUQt29Cr8mP57PCmkzVlsRr65lrmmd4KBUzBwslO7/oY7Hup/kyaT2DAinAm/9iO
+aWmHgtVelNbaDDGc3Jf0rlDrZi8D7cKcohTbPsLyJgyT4I4kRk4gEsfsPVZbaDS09B4eqw/u/Th
gHFsIZ2zjROgtpTrlBFV6pb5QUpmr25rSYZ3X5S9bV8C1gpn2ESbl4OE/d20DTW8almVf5ciBXA8
zRFCfWD4MBdlLsWBBhNB454BW2/mWivBJwFxgvfvqGXa0xxH2yGm7gzW5weSrAFN4if0mYw+QcHD
VLVQAQHB9rReNGcgwpHFD9GMmA8zGsGTLTViNUfnE6u9oYvAtUsWh3nOq6Nb9sy0rhZQ8REZ669r
0BOcIUuDbVovZfL7j44YftTULrtDF8kw37/X945vKaApCr8Gu75Xn5mrrG1ka+Q51lMdh9KHCdD/
yQpJxzW34oZ4aIyeP7P3dawkXQEZ08x1aA5MaG2frA8rRoRlG1FnDP66WXToBSPvJBope5nwyvYF
06ZHyEhyvC0unug5FcOmM5QIDp0cSN2onPxz2OASeo2+hoUQNSEiVKpqF27g06DoHeveq09UrS0v
jiJRwlya4lvThoQdFzwDdiaCKOhfW5yZ55NTsSQq153R40Pz54YgtRc6ule7curbhp7xMw/Y9pxT
JP4hXkNHGkLPIjhMJoTReks2kWLRg0jnQXEoBD5Ijp2wk1EBtqu1K3GVIc4osxaYYhtvl2j2R+Ap
GihyuxNA+26bA0E60SpIH7gda3UqObqX8PEoom8vLfIYvxDr/sZ3+PfWzUgq3pohaeEyODNtm9Qn
LEtpq2InSYKxijqIEMOD0dm39nGZxRuzsjzCD4Jnpohht9V8EHz8s771CORaK5Jtf17WvXgr/FrF
6qj02QfbdRjcVvM5FvOtLqcSNYLFErO/HC1B+YHpEFKiB0snuyq61TGtOrXY/8oPj1NRRQKRTllA
pCJce59vMwljZgr28xlkT6Moso9wqTmzNxWYUPBXY2H/sLWA00ThXDiTjiEvuQ3SrM1201eyErY9
IP385s+CCOY4GqyWWcYKIM25Tbw5f34s7nKpkjIYTiRXki6jM7RqYZvdcnWgwdHNqH4T9vCYvXM4
i9SCN+zZxiP9aFrFXKemFtYtyoIG6O6DllnQvS/cdJ3+hg6qHlRd+d42WVWtfCcE52fnYTBsrtIA
8RXx7mSEbreUBKZ+xM1xr3bOkmI3GTvM8fwxA62Min1MP6NaskmdfS9nK+fXnGPs8oz3eHEsERKT
NNzrNEUG+W9q2nlDL2mN0LSj67E1JfHY/8xbzwwwujGLqEVu93WX9G3U5z6uaJc6jiMpM/SHYSkQ
ACmktiiIZVq8kH2NLppTKd2t22nLbCJdfAmpYOTLSEzWx7YuNW91eEgCmNqmcYUsnb4Hx/06M47Q
fiirxhcCaTiO2/mmZsd2qv0HsOG2Jj7YPtfpp/jRFcVheQaWoRVy9Yp/MvmYtIbBatznTI1UIMB4
AdCmTL0qgcSTzl5XZ29tRNFD5b6m045PD+LZ1d+FQEiBmUrCnakW5BXaj/tdi/7gz2ZmXLcp5ell
6azew5wgtOq36JfO0Sp9eYzrCBVtjhG8w7si0A7OKFqDQdyP8riHKNeAO2LefJWILgT+kfCsFywR
1ZlncAG4Mh32iyLVl52uAZXCdMoq6xm/QvilWd/g5r8CYUid+burrBjyPKp/P6OanaHeI1qqxaj/
zmcvk25RPgJy0oNpgGYILGYqhXLehKbLwttBKu7t5giRm6kBToov9KJb9wlcMynKeiEZWxUJR3LW
Vu2FhKT4QFFq3j0qT5qMRgflfs+KpZ1n+4JMng7I6zwAc1tjDygfZFlUtdU1NrkhsGJrqOYNWiKW
bjWm6J+V28wANs9/x5Pz23Aa4iSel5d5RjlUNAFPuKaIU9F1zXYAmPbFaA/efxRM9fpx3fF5rh/N
rvXCd666cVTUqk+HSEWCo30H8rE97i9IFhFukXUUmJS4NKbl1z3msMjuP4KK14y/iFahnalwyFtn
uCiMjDoS3OyPpPN/AFMwMPLxDhCJpL71nXRMwQtcF6rguBxXbVWQLTir5tNIJmcoz7/Y2mp4/gQU
ZQQiuL6aftRj1hXvgHF8ax24ICUCR4SoMdZ69w1fvIm8TFDyLkRxaWycJYiwb/mJCzakYCI+NkqZ
SMd0ISbwZlK1hkcaaxNCfTPL9Dn3GZsNGN/eHpHTU9R3NJqczrP8WSEIWVDeBI+gTdlOKRbq0lHg
vo2DC4yQEGCkyya0LLDpqjszLv2l7fRiO9B/2rCR0ZwuraAUYf2ycihrb1Fib1sqgP7gqVZ0oPAr
Y85PQ5bI/B4ToB0DrBN4pGQiFglXuLjrjnNs0BWzlfOYmVaBaxq8DeTNTdN2F3NIwnHhASI/LirW
d1dE8JIaXB/mIEX5CWkon5Mko35l8kof1u++OESDmSxJG5B1UK55sQThosU3YBhvibyHAAvuu0cI
FWM0h0XydObKSfuZaFhnUkU7GuPnGcrRb+J85WSfDKv4PiESOfnJYTXuxxc1QSzy7CtTtC9u9swG
fI+XxrB6IHhj09ijVK3pE8kiijE/A24Rjr2X5LhxW5Q4fLk/m3dqcc9f2fsMD8LkVDq4YX4ylL3j
sLgs/BXCVQCxFoU9KFCqleLawWGvqVDquQjYIw0oR+Bxty2ZfU6BYhFg/myk67xjvsF3fhE7eWDy
zODsXfPw/dY0eXbGXxJ8Px5e2JGjF2i4Ovm2F+casq2mgukclwFtjpKirZvl4SoNbV7lAs4DxBQt
g9tMnxpEoXaJosILTo2RZGd6Sh7G21QoRx6U6Okefy4KDKFHR6qb5sHx7wP/qJLmLE3mmIhBAIoB
ttJZsfzBp0hov2fgHa+ZrHktaDbvhe5S8WOeP41BNsNi5B97EcrpvskIeWyFyXz+oL4kS8BSTyRS
aGnEcqWg4P3FBOsxEL5hkWLQdQAnrKs7CozxSDZx/BG6AvECV2qc7sBpL0cW0G5yLEjSY1Wm+us0
xpndG/Y7qQW69P6jCegDjysmpT/g5ElGF+mJjX2uUOl7Ysi29aZssU0E0XeKNv9EJ/YFkafiFvrn
CXf6YtaqtOUhD3LBC6eop/WDS4CZ0EQgWkwvUVfcRvengkxXhqvkyZY6xGdxgIkrKgkmOkeXEmKc
mh6NGnT8rjJ8BIs2oc435EcALZhub8XDLNZ6ngZkm9OEEgCrfxCTQnb2DaQ+sDJ7xdwHGpCQ9BAJ
8aGtRsZobDtdjqnxX7u//8PDQ2HkqKzzh3qxd8jxnDDph/3RI+tMFWBaR5FNHUwXgJukGHaRqseh
8LV7A4bMewcEYvw5YAY3/BwdVbjoeATtjih7rQfoCuwGfL35tmQQbDC+atVhfaPQh8pKjLlpQ4kg
fO/CEnsvxGQdosw8P3mp/mzgUvy2wbtFR7YVcRvEiTgc/dQUVJU8Q7dQolXZuki7k9DAdYA2gb5j
dCnKPYzn6BXDAK3lJLAc9ofNBI5MCW16lSyWes2LTXzV2/N5yNidA1UmCqphMZ/fBDjoVZd/14uH
LAT1cZUY4fBvy+MBerdQXRSOI6WKyagFVZdFIVx3XTqwb2nLjFKpInVi2uf+0ptrfqUDdUJK8Xay
MyKDLHrLjhWZomvHFRVzzNkjD01hjoYwLphs0Fo87PEWz/TUZ+6gLlLqWd3UZIu7JJV+QakwRhTv
WjBejzh9AwcvsuwH/RE/TKSIsLh6mMkzPfEFvxqZHXri4UenEeAMUpOBv76mGc2XE3IgiXWOXX3m
KElh1E19LYRcHqMdFso4LLIpfAvlyen2lI299Yuz5BowlYQdUlUcVl4lv4u5gotjfj3Lw3pJWkbN
IQhDccc0i9bUeddTL8sS8/SQb6KGF0lmvvtYxZi8HBh0uc5dnOeB07Swngb4PvtRShOh95xqDaqV
CDHyK/K/v9CkMpK0eRCK771du8gFfWlmX+iQkn0AG91GOKCs8hx3fEg7xcYepiERWXx/uA1/uLzV
xdhKCCH2PYyXSjrY1kfy17qNiYmkZu6YRXEFN+8DLmLD4mmyATbfDcudoyJ2ZBxatpb7p2k6BdnE
pOmcRGB+YEwRlY9WI3Zk1EPIXfQiLcxqo+BJ/qKC5KqYlzTJwS3KWV3ZBFV15l/+631xabB9sJpB
B2zYqwEDbL/YCKkCHEQ2M4xUlSUL6DS3ncZEKS0ZW+KO/jykbBtOLq5RvPjm2103pcRFavFlfZR6
kFO1vdC1r3GrWZXQc8zswg7XrHI4VSYHcl3xbao6vpucIHr4w5aTbBPpLM1sYC2a+uewLmnRenwr
7OQARJmeaL+pMUAXDA8BXvt1rFPJ1Uewp7XBf8tsiKoUgh4nficptJ38PLwJWNd9VAWNHjdsJ1lc
H+aBl5NVgVwdTDSKBtCFsAZhB4298HY+RgHJm7us7dYnoPvwLYlRthlYcQpmZuADS7j4rt6pFKu2
XqbidEOgznYlsDacCKoWo1fsEy/fq2809cBwajXfNkCRGu7NgHFkqlsqtx0vbDuwR7PLwb/0a0GY
7RNTziAIhxVKcPZTIK4x3tJ0ySYz6Uc2OaIfKnESysnfTQNvwzSNrO1T/jNF2qEKUYy++OUsQEUM
Nh6bJBgT6TQB16n2cnHWd1HEuwLnpDvNUUJuc6FgxHqiHBsl3YHTfzjNUbAHUo3d6DReczlKZCH3
6AWF1GDD730Ye9mxtzTCSkedFZct0ArRAG0wg8xAw1YUCCw0AzFjYGqkQHwbtrZUVPfYEX1m9WRu
DRTjwUZKhRcTyz9FRL4973pnNxUsbTro3CS0YjP6RtYjrlYiFF82JBTxniUyZAfMbXppkekLLJfL
dCQ9vWl1gQgWV1qut+oh64qy1RXwJ/lK///arzdnnYGQa3V8cJ84DJBba70ISeos8fz7dRdQ6h20
mlJvRZjuqmK4FkfAQn3Ru/w6XTe4tBDUkFqdDJv72RTkZ9T5ywq7gNWlulj+PfHK0WAjW+K1p1gx
RKznAHDFr+dl7TRibt5egkc5HJIi1Bhp8TQI4ZJ90Z5sc8D0xqrtzfwuzv47Oig/sMmmJI47MfGc
6SlHBKhHGfvx3g5Bo+iqmVMAHDlW5qnXdMrQgvKKGX/xcvqJmcvfI7z3weT/xAiiQatafGvm041X
ibxtL6zgU9HpqpFIj/4gW7QVkXNMMGqU34hDv2a19vjhfPTb09kfeDMXuiFUqmg/qcn4WS4Ic+L1
ftdQdxIOl5J/IuA3htxP8DYV3t2XBUwUsHES5DUjCk913tWq1MSt74JMUKFRl9MNdNpNVR8l2Xnx
+eF/c5wPCk35dLZ+642djWH3wnylIGvRKp50wIlXzUKU7I4cAReAHKuBmHusS8qY3vgj9fIrcZEl
aVnd0Q26qXYdFTazMY9W5GMKGjEoBRM4OW9YyPTPZANql9qGZ3Bm6/yOG2nHUuqPPpeYfxxfEOxo
osHarOLwId2eUIr9V+fA8uzoAxa9Ve1iPrJJNR32K5VF5Plqo3Bd9vreGLccKc75urUGbqNvv/Q4
9BFQH6dz8DypfpUAJVnDA+8J0We/ybNPm8zpcimJgqwgAQr0HUBjeeM6UQfw5WSY5HqN6+1EI709
FqmU/bshHmTCF50znFUH6ldeY4q9vr5r4hcynqy1BzueBfM39Sx1k/s49nlfSqaeXlhWh0zZeWq+
1KTGvAvkWGwTf/d0rdxJvdJfqUAxhowueY7Xy/HRSVfqDqK78Om3VXYygR5EI0UtucpddrpguO/H
eGXLn5+s2spXelhcqVrg8of2XAq0bN2U2Q/Vhgyoz2FVSpeAWIT/GYYxgb1f0W7yrJ3W6kI7BSk0
asSIbd31FycRJoo8D+20nBmgj6ILo51KaBfmpYls/h+8FRCsnQOu0tFWK/d+x9+U1Gv0Ro7/fDFQ
RoJwIyabuB2sYLlQgPos4IR+wplKeB6lgCmZm830Yw7fqId1RXPM+exBXwlAbWUOoq7xYeInZcqb
O1phsI7Sw9QRem0mhG3dT3tKBc5jgfAwpH/o+T34PkGpOjV1h8a5lVIz7j7RytbbNhm1ubmvlZCa
KmHiOj8E6kWpMeG8fwX2vJfs1kK1qv/xOe6Bv7rgBM/T2lce/aiqiNze40Ou3X8xs+Zijy49zDIq
RslVuTyHBClPEgquw7Qyk+EBYyZEU4oS1g2Rm7YOSiEyLbFQtzZ0qNpTbMLObUGpD75ZnJnvV/yQ
MttLYLyRW+WHgjORwLaMwXxAUEB3hqvT6iYFsrZOS09Xog1ENymbsLdZDnpWT7CSLN0ZrkxZsPuJ
1Mud7kWffTLzueO9u8xzPedn1rRKuWKdmjZitlLraVVo/HHRaX2HEsiiS8wva1Z5UFOfQDw4KRQo
ZxEpEUGn8PFp22bVvVDvaMmVEMrPSWXynmsBIWRXcq4PVntE3QqvwNtxcGsAZKUzxsKN2iQrcA06
Xc0vPyT1Ue0rW8uGtrGKtKR+Bz5kCXwwktsr9uFcmQDUasDtIvRLxAOk7OhCrKoFb94BRR8y29Gm
Nc5SxrMwKlrKTOxfD3a13Yi4j5ROaQ3l6pDCusxMntvYM8EpXb3wUcm2tws0BB74MG1QbShPdc8P
X5gnpLt7vZV98mT2gv+ZBQW7ziuf31gZc3tAWIbb1Uit6Vzw7xY2BF0SokOvJh0/2Bxy71WX7PID
WScvPPArlE0U87C3VtpDh42uUxB5TtizURyWNg1ctmxlmLLErQ/jsaIt21adtoFle/5/5bFxgkQ+
K1m9xIi8pZFju5FhD2vSmvP6OBaOlgRTXjpn0ZnuumSMnZR5wc9FzPbd3mjDP4TDf6pWJ0I3kl+E
Nw3Na+r1yonhyLxGNeXqibg3xNw1HlIomLXpw6huMqEgF4MQaC3bNMSEqOHPNYQz7tWWok+mB7Ld
0cW50fHMwFbxjmsQgvUmNgP20j9BZ9MYVc3Wz8gaEyKMgQLm0NFtB6KlBC+zGMUPDsUKHHpXAiJJ
NwDNHJWu0LuELwb+pMQXKdqw0jg97N5wggSxP1wQVoH1XS7cOffrnLBEBorXqJ1ivkSgHq32AZJK
2yGtxo0wd5v12bSIizdtVodPrplQOyQxsQPN7r9HtBn+H1J1ulfi3Utv0CfOvzoXaScMIeFZPLTO
dbANaHtIQigoB0ir3+e2h30khT8eiE+j2rOR8oreazETcJDZxjWbKzCR3Os2KI7Sew6qiRWSVw+c
8U9jJUbPedzhdajBbjZpqW1jrnLZ+ALErEkSYCDPR5SxBE++iQw/UcOsxJWcjKVQROi+erQ9cS8e
U8qINEVyQu+EhfP7TY5T9pzSE48mQZ+m2K0rDe7dzldG1bNFmd+/p+0kyoCqBQPVl6TrLwxdqkKH
+09rcCm9dGr1xTx5Od7bw6A+eCZrIaeLQ3K35sQuRvNpevZFMnjZISY30ymWIHKBYPIlq9pQgUvL
I+OMNyamnp2GdKaH7RlX5lWpE8vVw6e+UPP4OuDHQzbv/IOLYSZrIjxupo5Jw8bNtA5I0dlhHJrP
HxbxzWKxHD80emFGVnZjMNUe1bb/LKGDdTn58hap3oPJQgjQb3ygkCz9hkr4D39b+N5OEbJN5T0D
Qw3IskXHuv8Usoj6b6AHnQWNnwqswGaTpJ4Cbf7HH04Jw1A9r9E/SVsIFozj6rfw3Mhi4nmgbXxJ
gX1DyYfJ1CcAfRI7eR1VpwpE9v9vfuox33XaMhmcsGALnY40BAfnKlnpTLno8ijt7RCdfmwezdrf
N/+4RW6yT1G54YFFgXORv2CHTJBxrhW8ZngphQlFB4BBDHisJJMny2mryPkJPQ7MYCUWohszGzL5
eAXRvKSWLnP98IxbilLwBTEFx69dMhc4Xz4LFZI9bBB7nvjvq4aMIyTNR1Dgn7AJ1zQJz2HiJcAD
7PI72H5lXBk6qw7gunc5Srhhf4YyJh2KHfb1xirh38TkUI3qKbtB6YxS2joQZeVjVVYt+WZWcxrq
O2H6uW7btq6x21G6jyzhsT/JKCEkOVUPIF/8sZI0q4cvLQzZaLVurUSSxWUCrkcW8aq2HHxHrCPG
KguEyCmomaA0S1vQmh3qNQx67aOEPx/igHNl1FYEqgQDF5hqwnELg9Gv8GrlFeL50A+iZZmHHlGW
wZLUKI8s2S7kO3AQFJXoKNgQhntpCiDOd1MG0YPfxBLofSXzNDLAr19tRIujtCFKCfUHeEg3y3eX
78OUcl/5vmOpmIRSxUFTbb3mhJ4wjI4qHC4ZQRpHBBrf0Asqwd8G/rLXTvU6oVMqqpUkpb43lX8h
Bz3eRWnWcp5v9eVDhJcmKzud3LzuA0i726xXFo7vsJSFbUFZHw6Jyz3X1mvBPExBhTGTakAjkvez
sRDSkOh+EOE9e27VISKdovd5eIciN/mr8nku0KmMWJbiyry9A05dgMxOxXx3E7VobUkX921Uano8
bfNX1blmhN94HPie9WSuBboNzxzK3/x2jr2/4dahSjG9LvvnZ254zGiauUuxGPltbu9pEq13iQqL
PNyAGA+3KzjenmA9sz1fLog6JRF1J9vAU1BcKkCKCzyekJ4QaIMtTrRXcFjM+d2YMIkQ0q2kQxpM
2CxFfvUTx0QbNoW60qG7qSHV+u3DYBzDr8DZHLEdMfzU1xGnFf8tyybMWiuKCFbD398MJzNZ3dgk
SQD2H6+dR2974TsH6Yc3JT1iI6KR17114rFH+pHu0ux2/0IbqbtJxNhcIneBQfewCGKVkCbOkRA8
mk5U3URaWdAVgsPdqNfSIlx/6BPLfOcbdNc24y2iwWqbNZ52e1j+zsxMGzCd784SjJFwOyRQKZQS
bBPVuLvKrUPyf4f8bZ82YwoJ9JzJzvMk4t08zPoc+eBp78dbp/38Pp6fcKoj1iyigUzcZazTCUwk
IpknjAZ1MR16aXVNluquGUQSq5qFsnmKduVrzzncyG+05Fs29kgUmcC5frYpYb56B4xSDak1ZKHY
YQCQ3+c60CrL5wv8G4JJ9B0F3mYQOMS6ItcOcbgzgbfnNr5Auw4ABX0p773KQ3mhtnR3G7ZN0cu8
FI7geWi5mPCH1LYmz2aEIkgOPwAEhpGRRGsm9x274QLWhwKfSTUefwihPyyQ/mtAZ7/64+TOViQR
Tv37GnZ03xK9ToLbPou3o5YCH6VafOSdINsj1cVXg1eaoL+Z5L+gQutqH4lHRwm2HKO0tPGAbBRj
lUKf0XOK9HBsbDMGa5QGJD+vHVr5SGHG+DcIcG+bTMSchUY8vKQyLN+FoSQnb72NYDrqVTRks/kI
Njlno069jWG0F0SYxwgQQSnBPlVFRWc9uo4Y4nIUVaswevhYeb3H7XS94yl3PTt1tyAJBQWYCGEW
8uykLv/wBy55UV8XInivW2xkC0tXvF6v0BoHw67t4suXaoDjHaeYOqs0OBDo6KsRm2AhAGjTsYYX
XuiLMQ+oXW2jn0KUFH8I0JT+C18WBPhPy9aSjzCkowreeeEAhfehy2XBtQmzFpp68bDNN/kFI09m
u/5TCF1YssNn805/jweMHmTs775nAjI6iryJrVQJg/82HyMc2DmWzdDAYlkVVWxacOZstKhjNLAA
tAn0xHzQn6+uW5ZD+IjG0AyE7cThLdU75sdg6RtBqkcVEp19yphA+MDJ4JJ+4rD+DT913Y+t/q5W
ysBdMJjU0vRZjLcbZ3gppNGcix8tLib48ruSAJhmjz+v0h0X1Su5CIpBInEfUtbMoGcchMYF1DfI
JLeL4gutU0mdIIj80HaIFqDO5tThoyFIph+Lk2TAF/31IybXO/XqDNHl4ebtuKFBWjBiWv1RW/01
kNKZfJ4QTju0ZmjwL9FoXvqlU8/AJslprifuZdY7ap0it9bB9oMmolwo2bK9L2T4KVlBeQ5iHgrX
0o4YLYXQXIfVyOu57Kv2AaIZLA1p437YE/Yd8oN/OPfPX0yZRQQYBxqXArDrLP9R2PZ66fOvH5J9
lvKZGWmuut1Qc3LrZP/TuLjmxHMnwjTHrWDvK7gbUuoPEYe/rR6x3BvvXAy4cXaN5oQcMCNKliJv
boQ6VG0F8BgCPPU4dUN1xsC6JFbtAKI4nuRO34PRU2BquZnMYTrVPAc8Ew7F6IILCnGLIu/l03OZ
vj0V+UNe8bLokAukiS3ovO9Pk5dX2osauLivVWJvK1TPJ8khZMzi92MURm/e+mtkBIBLEgdEHQ9W
nQaJ6K0oj/QPUF6IaR6AIdspOe+6dSmAk+y+GcsoGWFHSfPDkKsiF3lZqpfgWd3SUgkD2yeOK/NS
TYIHzu+tKAWUgAPMHi7R5J4NPJ9fHaYJpgmRTUrZseWnrXRlKwM7z5qaqgfLZ8gK21fAkMwad/Tp
+EqolmOJdoxFxJCYJy1sDMV+DzFQM1wldx1X1Fu9XrnGgMVIoX0xBrNt20jYo00xtzkvjlhpTc3P
Fm36V4c8GqeGD+P9AlcaFzAfb9Oe59AfKeX0/TQ8eXWkm1cEu7r/B/fRydGnCBLSvN//8vip7vhk
Kg1fKYVsN7I4pK5SMDJ8/X7q/JF3jyzZ/VhSj6ihnCJxATnRP2UUgR07fLoJJhxz6+8Vh4z/K/Vl
5qTIht9LAl3kz+gAtJjYKZhGjTFrKWZyGwyy7tb2YezJsVvnd74vQ85jwIumUVYjunJ0K/DZNy+U
NC/DacwThojOo48E4FUOXuGGVDcMCovX4L+kliw+8UNOl8+SuF8ajRh45XHtLiTvPBf4sNjkzei1
dWJSJ/COBrn631OM7RVzV2qCNIkzdbsTGY8ltqLPUhvgNkpD0H25o0M6b/A/xjqHUQzPtTrd5k9F
wsvLQQy9lIXAZb27k6YlZ37fwGcUSr/FsONjK0r0M468BbjsOzEHDG4LjMJ6S9gU8lDcs89eN0uY
4xSuywIVrFbUP1PGa9ZmD0hlblUupM5/AeuiNva1nVuwN1VuJQgIY/yV0tHaWmyjX7WzzwCuUjvb
4e9KiO/nw8HU5nKmLsn3vDPMNd+O8OkzpryaVqH99SAqtmawjvssEQvWW76RB1KbTQy5uHEVEi4x
mT590hERGdboHdGDMklsdu0VWknBELn62aVhrrpwqCeSAzSY7uEXIq/5E2hqvp0r+6NJVNwmxFh4
CJ01xalzCrjegyowbuKIPGGnkt3VAEN/qCaI8sHemAv2To7qVkecPCOwPLKZCNEMC4b4F56nVLu/
iVXcbzPqbBnfFVoSCQ/++zCx5jt6LIKHlW5uEyMF09lD9TJsYo0u30qCN+syqYRjhAa2TiXyMw5R
h2YSpZfm6g5jC4/QL/IyBOKox/hGz/SdluwG/S0a4epEEA3TGFa/8dUjP4fQYvDLh3kTusrJMTl2
rSkPWlfpwS8WuUXosXDkamfrSGUEsvt3oztEgbEj8schPjAlyrkEXkFZfDHf1ipi5zrLtYRCuUiY
G2TqxHQu+T1bi+kuTm6E+o097LdqJzah2kWQyVTvIK5go/qO/UgItS1oMoUZFsrZT3vTPHwAt6rA
NBfCPfEgXKcoGwcmIqcQVsHSLtUwC7DhEUx+sP+VsmBjJptV7eMqaONQa8BckvaagfjbXEPvlfGV
n++xRbe8ttEvqF6NLLpyxFqFe0dvwq1SKmwU4PyRdp0//PKsx8Vkf1vAEoMfksSvgUPfNAuOm84m
xcKNl/JF3umwxNP5NGZraNi41kt6H6mTRZvKiDZAbwdRj7haGc7pl4c3MYr56zcLe8ETtyBBQ1Rc
e9QCse+naCyOxE9LI+iUzvu9t3H4IQyDnC8H2FdnGtBwW+Dm9QDIvcSVDeOgm/6DN3LyE1I9ENpE
n+Cmu+pA9/3iU0IJEwzxxUGTrfd7i65YK3jX84gtVSa+wQiCcMnpWRrD9vUXE3h5wWdB2zOP6V0I
m6MpkcCzNwMUmrHUREs6/1dS/JydWLF+oTSpwUuFB+/XxgrOxppqijVu1wJrFMRZShyjzvCVcSVy
PaostYfB4ltvg514Ik/eTMp0i49OVj68xLpCvdP2gRQs0wh7Qxxeb2UQWPfMcyQMVFcIUVmpAfxI
c/Ua9d19YxpBh19wYvXPDqyfCC4IWmfyF1sEBLZcwPjWGa9qHN7j9eIz4jddZ+w4COoIJTSGzcTH
8xmOW99vA/ny6f9w2nd18xzYuAk/2SQHT1FTHQ0wyRInmmulRhazdK+e3D+NxviCuRLP1Kq1rvZI
TnXC1QF1fDpI7447Crcc55nxj45GJpNBsQK4p7BPg0P3Cs9YKKYsfLDhCOVyW5NMPn8NR2TuMemJ
689tNA0DOlA5PwUJxl5S7pfq9rJuTblwB8GPoEAdxoLDECAlZpkJ9eb9iWlOOEVzN1MIdRVdBmx6
kiL7SNyvCqzDiRl4P7LQj09ilBvVlB+6JZzayiD04+PTouS7NzUKbct8K30QrlOr9CC+I8pdA35m
0TiFNfF4e5O0nqTHhJZ3o/rkwnizMu60jXINQo5iajusm2rUr+kKEE9/KwQK4yVRsTpulxvcC96W
veOUCgFiX9eBi9ELduG4sBK7DmEue8l6YIN9mJmnO4PHymYKo+81BNd9BA7xtsPQ9v3kIZ2XBBaC
pQj2jThABzV7m5jKAo/ztwgJwUOfesAF0aKcPbghCc+V5KY2ivnammG6KwhrxYvqbbw2HvXJinZl
5eLxybHSkVawUKF2DjfixClOerR+X9XfRIvJ5DE48Eu5AaQyFf4iKPvauGCObKWplKImVNxCdDJa
Zuf2yIkjNVLBmEPSpnmz21+QHWFZxSxVvmPKdPgYqi5yo2T7m15GEFANul26uSzHP3FXKLc2lWMk
5XWfcP72aF70qy8DurFg3sbrljFR8v2xRCkkx8lO+EXOGdE2LsF2npeQiwUTqB3ENm1omru2ErZx
hpgjWH6dQ2nLmF5lrj0dlqjknIrtXen7DzcCYsoSUWIKEF9EYmt2YmSs6TFRYxppqpcLLAUiWcOC
9O8dKeV2iL+b73rKBBKcOAFPmu9hFs7q7d9HwB586ETGTV433z/LmB9pcrMxRjqfZGHvR+zLfh1f
fV4aMdY/7DmIeWyehdNLS9f5/xtfjlM/e3HHWwz7Pp1lerE8PJyuiB7YlLYddToLHe70BSaE5dC9
D2Op2BRTwvqr5+vAvIZqJtZpiRcC5qWGSP2dlEZTMC8HPWaxB+x0yIkaflef0iKdblSVKmcXe9SH
OT9a9EjtYchzn8GJKIqdVq5FT6TTbr+GsA7iu/0gD/1zXtwR0+PLHxm6q25iFCz1MzyosCL+428W
Hn7IviRNsZSFDrZEj27npVueqA2vDtdQn7Opms1g5ZHjE85kKpvf9qLAlcuZMj37m1bjGOyDEuQu
oVoRMEu8QYKDmvc5DIQBIC6RveZThFXLwG60G77EIxEKDYikNnHP/TAfJ0/Dr8cfxJx4bZKLdxQt
VYJzmSEf54Cghkr782xhzYymQPow0Rov77N3hYToeCVQzs+ZlzhaiB/uMuTqdTo3n599PbDZl0/o
awIDvdUU/IZcJlfpiGluCdABnNKtl2bsbKdAd1E71ywbD2tFGq3Yka2aLzGrWw60NmTkX+Kkk29d
yu5waz3NT0hdzcik4gzzhDBL6R7gDnDKXLt2EkER4VzYjwT+SR1EKwElrR60nkn2o9YS9g21Y1m+
ced5eXYM2NBl/Kr7LySwqkrr/l6VC2RW6bOeN0tyMThizM6F+wqjq5mgQ5rwSQz0yJJREHDOnzBr
mNDwMJFcafg4sCXChwarWRVlgxJGpgy3cZ08V5L0pHvm2yhx3wEfz4Yt2aTViOmiEXP+nuIzClWH
jj46cEySy0Wcmkl3PjR+ZWWx/8tq1APCbyfxpUVkdg5XkkJJv/CinLLANrwwgLywWRpI9N8dSzVK
j7gGilkKz/Mk6gUsLvcge2cpb6fp+UGZOimwuqcKGy0EaLZCEHhnBj0nHsCwA/Qvr4aH8BAqls9m
kmXBhqQWNFEE1F21VkERuVMOVH2q/tAQgW/KTnP2ESnuA/nsMPK1fHe04ToXp53/oFwO3SwVnxjn
chWssn26nsWBQgchK3tPTW6ylbUXeoI3Sv/9IJk5GYVY+B684HWBAgffSLgJh8QpdTfM9gxCpWzR
XMaewH020w8/y+7nbomt4jKnLIRutyTkhUjAbYa5cTn09hZC1tPpezVXkb+Huj7rzTp9sHmOtz0s
xLPhtiQd92wYsbU/iZBQqRzCKnugnLS0qS9w/1rCYplWHgwdsu8nS/0YcxwDq3nvS0xjC86kc6L5
CJWRuriJzW9rmN+Gd7OUnC62B4FXEeTJFeQ7yYItSLQ16SOXTxMI/MYUT0DjLs7N63zDuqtm31cD
Jz3m4FiqT+WTX6pypGxusoSEalISP65AE1ZmjtYtJo9wUzMSonX6U9L69H2mWnTMDIaQqvkI18Gt
IEnRhAk1VDw7wWApD1pgoFz9pLLe0bPFoxMz1Sqy8zBGYaznx+TnppkAKekNUavP5FjShBUqlqRB
qQovFpYAHqTlpk5Qr0QYtXxEZolXz08pgHX70t0GXhtwD6TnSKtY3wBj1C7w4mX+QwO4WW5IoqhG
rgZDNp+W+Rag60/17v5PV/pFbqRdGJWwD8JFf+E4yssYAlCGShGORAjANM1bn2h6GwGrLVQyXpyG
zGhhMOZhVdVNK77oJyGS0/TEMTyj1gppypDlOPbjim79WwRD6hc02QQHzDgQoidDNbGTb+RFukIQ
Byp4+136ElVRebMAxw2IwhkYShDczjisoenbm7t/WhBAvpBmMVR60iRBYDCzzfPPijz1qGaivonr
5ivnq5KEScLrN2PBe8SUGznzLr0qhqhyIuJqF2J88CN8PXizHESCBAJ06TeY5V61FdVD7zM/aVUe
KAaaPr+Da92iIDnDNbNzu8n1eMDfQbrGEezFBtIT+GFKRoiP/1yp29ZLf8lPrxcPenen7eQORNvX
Sit1Il6Q6Es4kECdI6sQ5Az4dUT5W+5ZVwzn6YFBIuIJhsnPyqY1KnOUJGwvlg+iK3AvmiQWu0S5
LjNuaL8D9PFfLbMWOe6Z9aPXKlqo5tyycBUIgG+L8J1Mb3BVgYR+HLsLwPGc/39OQfHVriGPt+9d
wu5yi5Cm9GBMfZAioWxXC9WbwKVrpx8qZNKABjuSAX5u90/F0oBOfl94I7kL+S30g6YRijnOmzKv
ovoxK5YsUZANTL5Czu3DDV6bx5+7PfG5pLs/IvjEcNPflFcW9LcTPVu72BWIJZ/AU/QcZ7iYuHd0
9ZTvs/jpIaaEbTqlTBsrwxBZdP6QHUJ31qyPxgDylHhQyaqzweE0/wiHQ7yCINDSBnC0n/33bPyX
BTz98hQYETzfuw32rvuPfXvIoemTeJ6tDvp/SWPETnB2d3J1X61lNjiNiYYPQwVkA6DtzYUvKlTe
xgB1o2d+CWmAeDf8DU6hS6sJ4NPEihbyAcb8stAW2aySpfm7uCNBCRkrkKqWTd9t4rpd6G23CBtN
RUbeXOovOyXvmdqUSviC2vQ2R6HtGgdyd7OEMRlb9UdKZptKwKNLUfULqoTmbVrw3SYai6Zxsf66
rlPOWZCLj8kpXJDkV+GezD73gxFMRw7wQ5YNPuKeAMtvVUReIRtpV7W454HyWLnAr61/zdlpf+qJ
xWecwGep1oARWwnxia1FaFrYD7lt0jTe7DsB9JFdbxjxNAc7n0Gojnyg04T+tqS8p9BEDLtyYTrq
SUbctY1WO6j/xCIrkpMSOro0cfdgLM9+qLSc3SDqrNLgEPlsvFjL+TuF5ewvO7yKsJntzwyIk8gq
ckWYMMUMU0rn0GVdJ+L2tbhHEOJCzvoAI4yv8kTX3f90+JX2Cq8AZOFipfU0ZqypJiqtB5sSdGNM
We1nl5yRcANDYibgoTzvlaTFgYTZEi3wiDOfxSYQGqd0Q7L23c3+iLzUHfA+1/CrvBZ+MHgbt6Rs
R1KwNeYelatKN1GFc6tUZpsmaH8O5ITsbLK1lX+i81nxSYn+swDRdzNheHn7HFzlz26RWuRXuwpC
Bplt7dakPmDAGcWRS7SqeBIvtS1thpUWegWjd14ahE3lwEr/YbVpkjry9xmKAq8/ly2hUF5CNYXW
Bh2tvBUtMmpgvSATT7npuUYOPGb+Kj74WS0CZTE75ujz2TIpjZwycE12CqriXS4mfYMDYnR4QdDV
M3SfUshdjAvVbbQ0w8APKH+F6n9NClzog3V9cbdJcyYrJxTuY5Z0r9XaUWxKTD9t6ZSDrxfqtLY6
SaH4ll2NOdo5AGG6QuNjKB8RUGWUO1nEx59vbri1zc0fleBtJC2Hxfa4k+ns0nV7l5xTrwl2HiMl
cQiipCw97NUrZ78BsjDG5SMUTOKqpoaPklOqNt/sdyR1NMM3X3b7PMgHw8/H5goOj80hG6G4PEj5
R2qKqdflhQu8j0MNqm6OHCR28FiDDUhIEvxRpbvymTeOvdNsYXITMrJQAeiWg8HrsHZPlr/8Ke7c
/H7rr9ESC5l3DnZ17rEl0EKbpdrTQqF6z8foHRouwubDleiXIGabTatqGOBzBqoqGlfXME5clnal
V16IRfykGxJvNBw/OTvcN+pnMTzlTgamAmOjSd4nKNXYqtAGRJc9/RrsCR8BQVTfm75eMoF+5im1
6y2Cp7aIwdZ3cJgp//gJsk/eGryTmsgHLTiVT8371sRuwjncszL2J6c2A5jdzbWkNzJivFqLf3kH
HmymtxbxQOzx+rP8nZaN9k0liWs0WA0T133CmkiTp3OlIJXpx6hZB8gA/LC12RdtrJJxRc9Fql0q
bHfY8hwzQtQrqBsDsR2Pwpd44Whz5LoUYzrbgDmWFIKvFPkqSuAzokogvpQsXVyc8R/DbKx7P2mu
rbRwy3VH3ls7eCjUcYQcFHWYhfYLazgsyEBiLXvQOMXEgVpXuAlS2/JHG1deUDJleaJ485AfG+A5
vxT8+mBGMi4kCgkbruAIosYaX92+bDkNO5qqSd4L3gT2PsVvdQLti3Vq3LWK+0SLW66QBvaHFslY
GOzNQ/xEdrJt1sSlOl1vRf3bwEK065HHGW1lTiMT+tLhPv2dMYclv0Kj7z52KBKeds3QPPnlsjkR
fJdNeEiKZgRGAzz33g6PVV1LuyVCLZi1FIhbzjqEdJ85oL04sVHFBu1olVlLRR4Ed8McE8isWuuL
o5ygymX2cmI2XbnU2OHfS9necnpm+HejeB4iBJgtJLUX9lTHP/Kor5Mw+nmUt9EdBHb/3BQL+t9H
oUg48YF2iytvo+a1ZhU5/hM0Rv8huMYs6r1DL5yptccIbLFB+my+yEKay1u/FRFiHkBDB2IdjrGv
FtcAnV9nDr7DD/w/Ht7uDS3xkpME04yQ6jMcieSoIsVDc/wNUKgTgOrrrOnn7VtfnSXXo0HFO1LX
VIQun2ur9lZ81WwlAAeEl+9mVJJWvDRm5Nq+Pa1/po2Iulohqr6lavIM/iwrWG4navZMVW9rz2+O
oKi/A7dPQ6quYzdKS2wRkvYfXcTWOaHo2IlxPovVOhb7iJOAztNLdMTH+J3QsfUXWRvp6RjwCI11
vNFW2WGAL7t5uBnezFRThn8+EyHYdavOmuVLiOOeNmvmfBPv0525xjjbXvzuipvK1slQ+Xz+N/2H
zpW8ms+DwgPqzjkqVKCk7GK38K0n10OV8ayzEvDkCo4ZtagQGXhZRcLVooAeIvGcTW0xCHHfJ14H
boW6PC4oPFfGf4vkAN5lXT6jpaUTsyvAcDfRNA2V8dj3Tm9amN9EtrUBdnTcz6ASSLXvuwsFOqON
pqLTCFi2k1gjsHCXl9fDMfpMXkJFc2paAavny/UGrJIknkT5kV+aW+f1u91edBLUSOgAbu02OaLO
fd8sa/TPnvDHZiwlSjrvSIt+Usa1qCFxoy51zhogYmFQQo/Pyzbz0upKayVed5GzxnfemDi09ZM2
ft4gD4v6raEJasvzYZ/74PP+clbp1sKTzt+IE5wrRs6S26yJuYVE/rNGRF/49LWQUNeiuVFzv+ad
mFytk/fR1BenkqZ1IpQVQWCnD+5ObJd5oAyvXYD/OoF5GCH8IH4BskldXhG2cABP102+3ThWrY8Q
Fiqlma9YPwszA5yVVw+3hzgZRutu4OmUrsbmy5XhDNsgxJS1PuMjdaS+YCqLbjvTuu32ruO/o+a3
IheBLtpRquijIm2qOIVd2IUP1LmlWDajFCbifvRODIELDY6TxYPy0N8+SpTW9uVwbPi4xOOPvu5G
oEfSMDjbp7RIAri3oKWkPV9JCRdx1Uphz7hC1GMbsN80RO0nvppKvcTugYeV+d/mLHuT5h0L6Kyx
+RwenXHCfPKfIlBBri+Zcd8Opnk5kpj0nYGPVw48gADAcRNbiTyTPaHAFwVVlzdpuDbhgPexRtH1
h4MzWKkTnNodzfA5DbxFb+mGFSmIAs2MEcEHkwAAVQwS+WOZA9oUQNgZPUVPmwqXi1F5hjxfRlqv
CE9a5i7nd75+3t8VI8VQqgAFM5vkGVURnWOjpkjqBlEaJjJji8uTa9d8hgxE8Do1QCor8FhwdR4w
hE/DzcokhYIviyVvbmvd1vjCRCeDhaOITMYhbLCMlHTriLIWhfkokdRdiFF1mE/zHMaCuOw7qfWY
MkF4zILNA7GbF4/rZwNIffhMOQOsVB4B4yqqcHdrNIKOrF1lIoKRPGA1EAk1VZqR0evOwFK2pJVu
nPi0uG02ePnN0iiRewZc8W+PSTYpmJgRJAupy0XWy6xbsp7bybfSWoh8jpwOi9vqYDxNT3Il11dt
RPRzgT6D1b4/yDsRS7Q/r8UfCVzCu/YfMaN8W6UTtfIQF+pfdqdq0TnAOYu7Hy0JNtSyQdqm6Vk5
AUPW6uOSk14wavgPuk+CLc86WxlmgFEsYCHv7Js8wXgikM43ih6GgHzn9Bgvmw0ZE1XL/UgYKSCq
022NnZpeCj14QjzMTm1rfT68+reSAiv498x9v99Ay52bIW/AuP5Twh/196+9SRKaUGY3s1XXxHhS
MMdMygilhvhccdvQZohWyHiE3So6upbt+AH5bBs+addlDBZHWGkiVH9NJfB70HMH1Z4m+O5ez+bV
Sg7Xbjr0EVE9zHLaxf0cr2VMxEdr1SdsLxjlyVJ/eRijILV2fskD+xijI7XUhrK4JiSHWX1nfgcI
uSmxyOQVHx6aV8azCqaRWdSg71p6r92ejyj9HvanUszfmw7v8Nsn6TFF6iijT1G47VL2xMrc8YPM
ciJ7el3lU+fNvgbceN7wQ4DLmRXyzasWOVfv1JVxP3+N57Ige38B/NqYvtHFHSRfvavsItQLo3OI
VLTMgAsxSP7nrtR9tsspn+TBQUllN73uqmxfYgQugjPEXDUZabyJ80bcljIW/QvJb/GpatBWk0FW
si3LT+W2p4pkduSgjGKRFR3k/MgnO4iAOrOhw3AWo8yj65GWLbS2H8IACp4tSCvGJ7NCOBI/oP5J
+rApyLdJ/qUjoquxsHx8s3VG29VPmbEqeAkf55EQldG0ehSYOoi3gPBjYR6Lmi20VNu7FFwD6pQT
UsbuC09yZC/XG5Ho35xUjGTsjyzqAxSOdb4r2GRkAx4aaVvGQuwq7k4/1E2G9F3IvRic8+m9nOo3
q0p2vSLIP+HLIdbKZsWHVBdjc5HZ0whnbxNDcPXieEvSRa3UTyLH/PQBraTFe7M4zqZgv+DVdMqU
5cc39saHU7OOfyvhK/E92nOz03IgY/GiDHRD5ZqPj+WhJT4sygrguQ9mq7TWeL3ghleq6cMBHACk
fctEwQuhkVlN9/xzSkA2GH3jU3a15KdLTPNFpmNh+QEt93IPG7q6+B7gPnRXAnRdYseB+LGD1k+R
jpGPe4ZWE5k7jXNdMorU6ZADOuP6lG+H7o6jbDsoDG0KYuD2IaZ9PBvdZD+gSJ7/ynDaefPb3un+
hmEBNPCIGkurb/OGzib6ITwM4a7CdjlKACIYAEaT98ei5MxKUIlfDiZAMOouvEnq2uidzjZJZLGf
kM+DPicyx4bhcXkFir79Tx+Jww0IZ+5snu/SGOjlMsBJ83Acu1mSU90JHwUlO4INxorYaf5EBAPQ
FNGU6ZudUCI/58gwXqSYqB1dEfAtljDZ44JdQ2blckvmIxkQ2fnCzvU2AErlwBr0/8oitfd51U4B
gR6gM0fbvXJfbVvM5TPgROROGAdrb201apIMtWpYn75UdsBJlpmpl5y3rzifHspbDqyXN77WwLR8
Dfc/0Ehs8+ChmYdy7jKV6H/bjiJTaW1Ky4odGWA79lTQbjeH4IzM3a8m/lsD5AvDrpd6WlGCQ8ZF
y8jjnzGRCyiiSdVNTzE0SwL6YzuEPpt38Pc/fiuguzyuwAGarVOSfiuLuelAFC6iwh0xRTSSQ2Eg
Yx4MlIJDYXeGUC5P1FIV4spzsaYVgs6o97enpsL2ZWBuTunJS2PVpQwX3chYjqhpNRKb66jzlUqF
wD8fjc9JKWyM6BM1KJ09RafLBykK0jTmAMX1AD60Q4T9Hbi5zyUa60J6t9x+TERHwh3CxBU8LNZI
ETUO0uTzr4yvQayKsI+/TGF2mfZXHxJpviaQegJ8hUepQ/qLLByvW1R6QkjoTi3H1+JgyKDOlxFP
cal0v9ZOZ0xLp/YXu6xc5w67zsfPrCjT55oll+HXWSa80xAA4fty0WRTQV+4qfd1L50Z7dijLC+H
7wGF1aHSnBsYYAosJrJJrz+6UyodM37Apyx7a0gDi39v/nK8PkmjvSBl5idJohBo8Ygn2X9gopte
uPTm5foosV/IThEx+vCo4cXlBjlb0Vt+949Lyu67phHbW6XJ/71mfpqliqzQ3OWFn7o1rTAnpIfI
Y3cGbgeRpH33SDGRS8mEewtEGl6pXrVWB3wqqeQrrucvenoLFMuJVYHz35jQ5IGFv37AQ3xfWxDK
6/Z6cSlbT70qvuDULXCSZwFraGP6aGC9qOc/mPqtA0UI3u4NSDOSK70fUiewX0t/dpGfazVNrKWF
+8oxilnqlN9Og78xPLmmQmKXNRT//TpC+fmsKfOa44VoVA6Ux37KHkCXv+fcUZfjJQY7PVVtCNwk
jc6zk826yZ1Ntm0512d9vfilUBwSMBTiXLbRBApINFYo0hfunTG3iiwwmZDlgwL6Ki/a/S4tnJYC
jg76wjnfZ4WY6KdCbA/RIMLA9C4fXWs+mxfq4+RFBgglRya5hricI8NipiY8BdfNcmujBdT/WmyH
aA1MwbnM5aNTQioz8wjOzj38nA+z7gv7pXbbIWfegphv3YDdFb/9jvT758Cw3ZOdtHmkE5r0Aebk
7rgy75wo6EcyiUOdu3tcyVv4066w3T15ZPxk6T7c9L+Z4GEDIRbT2DxtLkGHeVXrsgFCmChAlVhh
1/ih0MdtDMGCkr/5LnFxuUaNkLUk0wbi0Xc9BBV4QFLd2+wBwlhSw9QE+WzQJNChCrNEaJMs2CNW
bndcGbiD6T31XoHYYsF5OUgNQtAnbNrN/dgqz+iF3RmFPD8Fr39oS4uciqj0zPw65nstUQSjkLxh
xZuZkMASfr2bxutbmu28xS6F/qAtKsPMba2GRifEIoCYJLuXuTq3RDLsHQJCw1GW3k81Ccp7UY8x
bitNBgs3G6jKdAe9KDJWnr81sUK4y8JmWbd7McjRm+dZLOM9zEZ1VYXqMNOTP+WBNvzpiGIXgOFy
+7NDoK/vrVmu5bCSxQmvD1V37keOZNfpMgLIt4qfWly7SMU3yVmdvFKkFtbTcT+jt57TMsfJSi7Q
IUqAJMycZDSWz+Qvo3eFbz8Ex5eMAn1dLWvg0s8XC3wpA0z1bOyl5lU5fg2mDD7SVGEB6Z/dU/n7
yzERTGFSnNlXmTIdE/q8KkyHSopNfasMpmWmGvl8BQVi6pBX8Ed4gVRAYNiwq/8FSOZOyfDrqnbO
P2fLDwVStsbS0jXdIVJ42GGbIjdcGQOr3+X4PZ2Vr32iAzPoJ2ll1GR9Xl2CwZjbTbZoKnbsFkEX
jbw8x8W/YgW9CVIFGyTeP5Lk3h8fzOtVt40r2vRCrC93QkaQW0ZqH2UHtqRLU7+b6jr9Pc+E9eW/
7jILQaxdd8lCWy1eicVurzshHKZ53xZRNfdhNCIdBm2ulsTBl4W+HjO6f9vBOMrlz8JCjN1BG0Gm
JPCKbbB8IkfKdUZHTb56zmAJ53eWW8a5+mTsjNItfVghY5aTORTSVpTne4U5rnggHkSqbb0Tugvx
hCp8wkgrST5HWqSo7Z6BWon8VdxlRL8K0N1/HRtkRjwZM97txd0BM3Nv4dskaGAdF1nVhykvSHXr
rVjvUrRPg2u0NTceJX0UAW4+K6X1oyLpgPDOqY0/mxdhH6h2WJgSzpHs4fJYDJ8XsGcOdWObYdX1
RGRWkqsJmj58nt4K9czKCtjHkm9ndY7xSjqWtZKebnvny/56Rast9jSPKGiH3CR9TtIUnrUADgCO
FVP0TfO5hxT+336N7u1kpSlHrwGiC+wwHf+aWdO/sHkskEemVdx3tRCZCs+mrWeSGsME2FBLIQFM
1C8sbXjhebptpkvKAR+7Gp0tgBpqo2IMbKpF2EPiSKpR7hfacYuJMnyjhws+6/HyL3/hGIbHhUZF
TNGIyBCgWj9BsSyPkVF2rXQNa4GLfUmEGT++eMlehEYKIkYLqohv23C3VONhKXbp2LXmwjUFkGhf
yzPVExOokya9BbOhQN4iiH9ei4KXIe+VctJPRbsa0RjWR12Mpj8vER6OSidDwHDyAJdJux+0QxqN
BZH35dshpx0XKSqy0rxnVsMUHXCgDDL/+D1j/6i0HEYzwjBuGAkqmKijxQyyQyOwzcqPuETXRoKG
7gsnzod1vT0y95yus2hy3tViRVDH+PWaTbDYMJTDCDV5bZO9bHQeP1OWGyaprgrKAzJ14ENQm7W7
L2QMVx0mFJVX1BnrF8zBBmo5GKij+6bbOFH1zARMpykcABfODvaQ6DZsSAQsuR+M+m8NDdfDwnPm
nxH4XO6i+RSHRNGS4r2sI/vKMppbfSDNhyaStWOvZe23Z8HFNg3mng0cN7Vkbniek9uxNydh5+bA
fRrndpbuFguzssQ09ijri7ar34eNWgVa8QbgOtK+DVynHWCGbYntwFeJzDULAnNXYj6jmn7XQqd8
ucAsLRHJ+9kI0PlzgvXi59C9uxTOrZ5tT/F3RoVYKQ3NzbUsxD8zsmPGhCsen321fuMybyVa02St
IKIZKErZih9Z+jY8bdKsDNThkLPYYlxoXEuaPrhDy+3nr+RraIqIOLwRzOd6IOh0tssUZaXZSVgN
CQZlE73AAQQk6zRuYPcT+hNdSlj427jvkryh4F2KpBHEGIK9O7s22otO6FRzKxZGjIjzZeS0EcDv
EpvQCEv6V8Bp+1nOI6mZ7687FAS/IXAsy2nutTAdMq1q4WqW90ehzeMUSKT/O0p8nHp38+wDib0l
SFWUVw3akHcp+ZfH/05agrIWzSG5QbPtCemi/oVk3icF9/R+LPLcKox3GjRh/dzX4WHj5V9PnJQx
Doz0C/iW552bUzKp+6klISNgJXAQx5CcJeUA01GzcwtOMp8j3yzRKtQKzON2yEwLEI/s03aS9dK2
FDbrO7j2fstiFmN5lQT6lAQG8I4KA4lToesp8Cspz3XVBR/E5rDO3f/2PAw4qUVsXitfueKtdfmq
V2hVVRcTjGgLppY0Nziwd5jc6/+jliGGC4TWMtOzGQcPnmsuf7ALWuNBlbAqXJcqTTZTsVvPwZEW
fMC6q575qktSRhDNfyoP3lsdx1LWm+voLo+3dFv78l8Zbd8diYoA7Y4skzX0uEqpg5Ye2KsShL8w
xCHhu+tkmVyVkYP9s+9feYH/htKDEzRs3SsVkI/Q1yHjQFJariNC9ZM9vOkJPiqxbz9Wx1QuorIu
Ut7omYBxDpe35bilaUHWXt8YLi1DsDa/I4FDHjys+qSOSRVU5FKBZCz4TN2427+TMWKoV6rrdIql
3cMPkovhPTWU3Mlj9rg8DjGhrwMC8wvIxztJfm25j6MDaJT/WYOIKNTffPg+1NAxeg5d41bva+Z9
flcuMJ5RgplBw7c3CciGupKw1zmNjjsuJg7Qus0UtJUoR1GQE9betsTIh7qlZZE5r8unmk2BbYp1
DOWwHep+3BFlPEDhUkZpx133kazCqAfeoLqnP8LJmLOlYGMp0vFEvDVXmSDv8lu7i4974yRp9cnK
rO4oBm4/4utvui0nb3TEKtJNz3swOyQaWRdRmUHx/eTgNk0zPTThKZic+BwtJ03jelG4ou9Eazj8
qCw9oa8SBnyxEkyU4x6kNYoI7alhTFxW4BzxBrJfT4dFAoGYUEhq/+JM+PrY2fyw8iNyrR4mZmxc
wqpyDng63Wc5CPjMllkPaI0xw3WYDh9+9K9mNr8Qtpb4dU1lVWGjbrYxYFq9rCVCyGlZO4ShrDdn
dBB6QQMhM3GTX3lBiy4gsEoLD0hMmnj7w67GMBfOjzOWRGSEwkGvFTe1pWAIhKraCQ2LZS8cR8Nj
wmPJrz0TkqCLVpX42Tycii7KxvpvnTD0RL0LAcBSmDJHEYmBWz0M0XM3mw1BstLZDbfP1ZYFlvlT
J/l4AsUMWWKT9EAik5R7PCBRyMUlhExXXcnfpbktCFx7zpXTKUGuiDYjdk9ZMTVpgHbA921CuNDz
MTvdFks1fJiFR4L5EuFuBr8dV6aB8Bp7zbEdYoTJYJYojrprZZhdV436AORkSlVyqtybF5e0Tkzk
z1uiQf/BIGlwYE5O6lPQGtauuzVpv2g6CywV0OFBXTzG0t2hOzU//IFNwh0//X0zauMqCoPan8WS
3XNAKcJlJqgqAsB5TofzqIu8XI3AnaoJXpJhS7egjksqd3Xczbmw4kW/nMTmU/um/qexIdN/6WuE
w2us6E6e4dQpBNv1AOTBfBqYii6UxGt75fz+XE/AA0gwNZ0y4zGv4bb83k9NjXsCPvbiNHAFJLqn
u0M3MBX/6vIyYxVMPhx9wMp4aQaEGByutD3ik7HlaNQiDysVlyX7KbjM8iqN6C7T+tRpZ2ix6xwg
9Zot8fRKZv6Rd1xQ4FW6pBbGiKjBmhWHov0hIZNnJXaU8XrFhfWgeGvzdX5IIobdDh6RThY+mPtG
UnRC2KvSZ11/gRj1A4B829lLSSH+K8yy/ecMtIezlKQH6yno9kgnp79mofqTadI0qrXgdeam7ETv
DL8JUNXV7VFvbwyjyHBiTja27J0vKpxGtqaURqjyuueEajtRWfOvx7VBuVlbKL27yyxxArRaG8ys
YIwlk2XgLTS+2BzTkECF5ZhBNTctKMpJK3zj7RqnAZykdOSkwI8+yMAI1kDk6Z7mQtK+C1ps2+7d
keeU5jOCQLGeTueSmL273T6yFNtEXniEa+f56CEk7dcm5PHmM19JRaFigDX3KQYulx8pLvjZTrbb
l0bsstC2azPMaTuAELUgn9+COIcFuVH4j/cwxnGw5vjMrRU/7PljeTi65wGpXSmeXbW5Wp2gAChJ
ZijcVIzWWaZ6MMosyVzfgCqIEBREaFxrw10y3xMziJiv0rvolWjgPIlk81t8dukusHki80RoizT8
mn9tYRP4bVtBK+8lXd4StIB55AfbBrNKkRWmD0QKoDGw52+8bfvrLQZssSOrEDI39j9Qx+NIc/qZ
a1Lts6l11imTPuvGzrqpM0jcUUT5Ak59AvXI8kape0SUAwA7OO7hAUXo1inPhiX68x1H9dEKYxb1
4wfhCi9RP/NOkcqOfCS1MoGIpkByFTlYgSWuZ7HnjACcW8lBvAFVJwnJy0WHmhxe7fXlT2472zls
HBqB3V35sS/aSV3zuSjClMQ+H01GSCRx/OuXXTOvio9muoAXH6L118ebOgd4Aj4r6S3dMv0NE4Vb
B2I73+P9VXtA21M90pNzhv0i4QkoVjuQhL2J8zaWW/TlWC1qVHonuQJr0wcFE2bSAkXSE6JjPvM6
nO3WX9fbv7F629VoR7/vy/AOG5q5zcGjLW6eiJ2JazUEXv8S7MsEWB6GI0Ae9CVh3yS7Xxd6YIq3
ui9c1o2qw/fa8S9Dd9h8Yc5G7QGvKFbsl84cYXXhnEzgn4wXsl99GVqkHLYo+XP/+1R8F84wtSWA
rScVTaXFdWJpL7lr0iaKMISvHNCgBnCMsHoxasfqImKP2vWJOE6jujPOdkqH5Q9ESo8Vt/MPGwSd
ClJIP/rz+iZNS04+Nzck5HuetQRDWDrW0+gpojbqaKAbfVjESi7Yv5WEWi8RTvvLFzf0dOLmIDrs
XGl+DMai3uFBKcBJKknhP0xRuUJPrA0hOGnrGa1LGl9EsSaWwcnhsxQidstP9QzacjerL+UBSLj8
/EVsvN1BciiNxAfluNPfwGUxH/cNL1AWTfC5bn9Ewc1smSGXiPuThniIIXtAH8R7EucgcDPYoxcP
N3Zez8cXWPog8/UOi6rTHJ9LaCP3QL3ojn5EbnCZrqUAn/U+XaAPCMg4jkhbFP/UpaI5Eyaoyqff
8755Ts45B8YYCVhXl6hgsUvNAfBug2vq1be7SNiP+DVjFQF6sINv05Gca2dHGwdjCdwTBmoNz8T9
NgQA4KU+6qYo9zr4y6n0yhe0EQRpG4P/SAkU5QNkoscnLtz+kOi5xFxy92wyHHQoQTYLSIx5H6D3
KmRBlsRxJAxBBKp+zyLKlaurHEDxcCAlXzXFFWSuO4Vk7tbiUasMaQ4rDLKp5HkzbA0jrG5wrUDZ
pnNW2Fv48QOprpk/51zL4GLRVCm92UWv/BUoFyjNOoqJmWlbolClXxdLbtzEP78IlS9pPSWkJOJ7
fRKm4d3L+TAAYrG414AHGmQD0jrJ/b6Lf1EIp2uLr+uZta7tmBgzVpGzBnD6CD7MXdcpn5knIDG0
nqnlfgKf0ehu9QAoBylA01Glen+aLKlXqSoNh2xLlifDy+zQcfBHoOJgc1NhDYJrv2qdJT4c/OL4
y61ekCAC1oShJSadncKRQzlvlpNoi/4JNgYGdf9LqlUoWL9TP5HtPUwHici4S10xSB0tqey5b8t5
DXNgVRUzm3NEeqJ4Zzhw0J09wGv8Am5b8QzXHidTuuDbTX6L59gZrX5/cZUp6Zv8hP6XAjzJVffi
OF4JmCtpoVdpGaZVVGWc0OeXY8wvwjeYJYylmiuwPFpKpeX3EzJ41Cd06jXQthu+DI0qcY3t5XT9
ktACKwOPH37Sc9JQVWj8ArnDCMGLJe/kG/u2zdRvWsoufGKYzauAU0rtZSx/qgKTw60WMRPJ2cpe
AZV1lgQOJ/7PxkVy9IWcIKFAO+Un9YXqW/tjkatxaUOiPGXNB4h5KiTkuELVIAMxq8EgGV040wWX
VqrDGFUqwEqO6IazTUkuTfA+aKhtuJsaS4sO2pdn+ZoXWZvRZWH/1uU25T37JJ6h7t1zAdFDZXOp
tCw9sy00C0YvvdPo0zWNFY2UbRatYri87oNryU+V+GdDTadT9u48jp1Rc7kB/4vQ67SGC6KiHB5A
cdG9LiZ4YxL+F2xf8Gpr61O0LUqbi+2Gtt0grZeiA4o0JUm+j1hoYUKzzwoIRgawkWyMPvNgjgC9
quwYjxiB2zZxdmwcprg7jShgeE/sUNK50DLpwsiIVUIaA7WdP0wMnQ+2vgjhPWs9Ct9c3+N0833A
ic1Jff/AD2Lk4Gev3GfN3jsQdHynhYoS17XIKjChMJPS7KRy3DQN1qq6fL5kFFRd6aP7QcVrds0N
sEBCRqFSd5jzaGcmeOQcfolpvwwFIOLG2crccFmC8f4QLucxF8U+AOcfaZ3qrV4w3Vk0aiW+jgAI
WFXM6YHH+YX6QUD0CFDQgqfmSfKQadP8pjvue4XWOtD5LT2nL3VgKvA8IlZN5hglLHuzvATriI20
7YnOefNrlGMuyNfWq/y+JbFUqvhVgygwCgWH6JQnnKCYx90C+/JRLq8VXF7pffMVPod1CcrJFujM
HMxJRr88x8jdS1nuClTPnMiRBZRUbA+9YEffL2sHC+7n9dIr4Bx8Gbpfw0bjSPYn3YsnnswArUZS
lDqQktcvKrAdOiKBRliMw5j87MQtzAU/tiQyl3zTjhxhpx7KtgRiXdFJ2u3ZR9Z7pGYMq6i2/RPF
4a1VOctrEHn6MhdRHVESmKXaP/QqDH2H7FNmCSsVNe2GOVI4fOb6jyP9TdH6dDZfA4OyZ0EMJAg/
NBvtFnMptyvpEv+aLztx9kJ7B+zKNajQ98wvOlzOx3jGgmUGC08/s0852/9rGW99L2B+Xa3D5GSt
jnNhfVOhH9E+vz96KP1QRQBWl4HcB8RdefG4hnHyRmqncjaHfnKhH6d0Dnbg0/l7cYAiIvcribP6
Z9C0XyfqefvcoM6TSnBZKdGGrfWhtfj4nSMApk420jFgU2tGZFSQ4zPVqek0w96cNHLder+2kxGM
vWGR1FxSONQnSf3nasNmcPajctrVIl6dnqW4xHa0BeTzrz7DBfw54ylZaKbQbH/YkdlPDx/zbSHa
1DGNQUmXzAYUrktvVAtIHzKPc8RqnhUGRiiScjrL+nZYYpIAlYpxCWe8oj0wFHWfCcJdvIQon6Ve
U/R4CJL4L59Qh8C+HZrlmyGwjuPI8USwXjMK9/03C69QlqmpUxj0SG9s9UpD+vp9vzij8/eMkxCE
Y8qdKBO+7D9nQRi0uv574PDsAZJZLp9Lk7GZYQULuSicDpx+dk2PEHq+pNM+dlJT96+9Vci0XDRA
w2artLDseYzbvfsZ5GUGj+OfxpvFIRs6rBCGadeX5c/eGvU9RtAlOcPCuQpgd0KBbkhWqTtMEI/H
p+NWBeyPL0RFsAxdQtZcOd+d1vQbVG40fXO7hL1wXB0FPUe3B/+zD3r0Sf/czsVa4qPfM8nEo2Fa
jKVKI6o5dKaAEV35q396zkMxrmLZTCLXJ8kxQa1ekzTEYWzxdewQ1U50yAW1VCLkkHXKc0jkUNCA
GHEI17MEo2HQTeihtq1bdcUsVOiQ/Cmyl8DMlp2WILVwJ8MsUfHyU0Vy/uAbq3xlWNc75WSmgDcx
nXDjmr9Q+r/f+EtioBB0pBCj7ZG7N+5KGvdpquF5LVpDb+3gn9PJtYWxROEiFjtz6tULUxSktMxn
ojyOsMkIIiZhrmxMUK44zbyVc/sDFk5qFLlGB0emVKh/B5G6avoeD0YnQmIkRszMi2nnMmhhGQ86
U2W89Mxtw9K+iXCpIQmPTuLWHaxqFaL2NJupS6F+6t5+HULh9c4iLHYDfd+0CKD9Af2m6Y/FfRjt
cNJEECYPLgqR0R98rq55NPdHreIJIp5Zmu602rDZb680ZG8qSfoipAWOK1izHYf4OlC0mjrqmSTt
YtecKhkjBttNEnze0/6dOrdUj6jywt/KJ/NYlx0wd7JOA45Dw39n35t1pHYiKQopPw3kMUValpY2
pS7T3eEaPcdVfNWOhWPWhxFz0vfsKZ4sfWml9w0IBOBfbR5FW8t8SKD5DsNcxVe7OeXSSp26G+Mh
E0FDvfBNLnozVtyp2NdTVn2ItgRQTuB3gNZ3mG0pfM+dcYNMREkWjysruAl8Fy5OrOSLdkc7MD+3
hClw+3LFm4Vl/sBoJPPSh7knKfRSPmdawpnHgvuyj6EU8AbisREaOWCH1A5QEAOqZYAe4ai/XCfO
KvWWm1EBdwhOh8YdDbgvv9XojzT1uuXWXrASD6Y2qhWXPFmwMiNDEwsyoNH6hdOX0HFsw49CSF5l
5kZOzubQkPFFnFJ62aKSh3//ZS00pCr8FCtu8Aj9l4yiZJtKesJe4oS7TzhNMw26FyO/TS7LLIvx
3qtzsVdX7SeGMvRwRgVlxQ3O4Gf9MgyJwie5Cwrw0gGaLJCBHBuWAhGYKxe7eOqnAuUf0ru05JNA
4EPwU/leejHPddroyqVdqmN6rr/0GtFL1Doh9xMOIMcFPyuYYspwPRHs12AW9WAtFm/02t2VBJdf
ZmyYRzFIrN3vR7syFBky0lRPrFWiyVoKtk+tJaNxUTJjD07ylTJPXXu9gNbqWJkbyP37wY1SC0Wv
AS3Mm3Ns6liwP8n/lrsGIWPfq4b5mImV2nPCGyb4iinCgF86zlSHwTIOnlFjs8aFNeggoG0MK83r
eU0ePIpvdiNOhgkxdGPA8YsGFJlpu75xO59KhzwwwFDfc8PnuWGbIMigACHRxI8FC/Z1sLjlwG9p
YGqXhGO2YrvOgBXBhh0E+nGBluckWSSB+izB2hwkev21tlkO16XwLp3gwq4lJuJ0a9O2F6Hpy3cs
HeQt2+Nww+2sCne5vybZ4g/GZV9TNjkt5c2FixdePnjtzzfFEyqbKZsBH8MgeuyuVrmdNEg+NeVR
uRdM2/fce/6HuySQL7+BWHNZuqTCL9a7Av+skvStU/1ziSceahIyUKKERSVJSuytwdUHShULCgeU
vNDMl833l9KoE5izqlaiFbs4VkChsU5tOmiBGOyEHbxCgWVShX3mbt8MXSGdgXAq49AzgLBRoH2j
faA9arJwBd9x8rX0ErESg1cloyzCn0pROsfC6HHbtcDLWDcnira4r2vyqyGN9yY+T+IT/dbiX6MT
11Oy029/78pAgDgc2hxUn1M6kNLhBkXspm493hO3FnD3YkXco8fsZhKeYeZevpTYyNkyNJydJDzD
HQg4FSnJ498uSPAY9KujPyYvLgxQCPDSIAIGEQ9OVq3NKEmJeZHNhJL9EKZJjYp8bFQM3GOqiewA
Tk5ksJjDUbK6iXP3rl4Ah26XStZAhPXSjnVUJpNmVkcgJkIiA/ba74+t1qih+1+h4jbL+hkzoUe+
xNvv8eClMEEhmf3eieoNt5ZFXS7xWkGwH9L/jpRmydoeLkXiVFfyYW+J1b/Z3qI+Rr2lo6BbiWmA
JVWo+6jgZgbXDySDqsrBB+tBKP9eZ19Veb37UCX8YA4Pqrl45XGf8Tj2Uv1pkJ7ZPsu3XFQuQoeI
iw/99wpRpY6MfzNIZfvukex0e1QT5ck1tZRY+wn1nNPvSPwwRQuSljZN/RIK7Gw4JZqe04dwHt3v
3h012uWu7A7lz1Da7E+IsfPf0IXq24CytFalvSGH++tWLIvJ+lV6RcYlii9KnrrNcrFcZuGZZKW8
t8/YMBDdn/WSQUdHC5mszGYMagCUZBRHZUDush5fvb6SlVaYTiEz8ezzQj6E5LOWi4RUBqfnuh5U
eibhkfBN2ra7WJ3EgEh7HmdMwCurEe/HaH69hIF3tjEJ7eEEex5prOReQQXuhyZ/5HojXVlUloMp
QBWi7y6PYQDfUUbYr33IOhkUKv9rfg4ERZhgMfHRs4wTKJSgx+/CCMeRpto8qsnXYCBnbATsk8hz
etIBEPKAXoL8Fm7X9vxjFyskelOiM9Duo9WcbjBBXFJ7WCzSqL3eCT/bfJdqwcLYsvECVQDcPW2w
TtHmt9/KqqoupdI59vaziyEt8MT3uJ9XVExh7I/x3IBDYUmGCz7ePisSur4m/aPFCACl0QhFQXy4
Qp+4L4BLjjMG3t+AQCnEcv3ySfYGDnU81SMZbop3XiGpBtX9rm+DqB6+fZfaXlG9bOOaH5PL3YPB
ArxoS4B19FyjL4oC2MXns2nlW62BHrjcKEJxR9/JJfjDe8D+v4ky5m28mGA3/5q05sF+DlJeG4HA
C6pPsmgGGsFYFd7suabSPnlUT4VrUR0b5U+HrecMYdipn25Uoq57KoZlD5FKZAfqeOQXlZs7hYBU
rpEoregk5v5WviA3Y9KGLcwyQK9fIoIHCW4nxZk9oF5wRwmLi0l6puJ42aTxzOnou/0agDl/7vxy
UQ7CcSgpXJYGW47/izkX1oKa+g5DbG7Jj+jHakwdsSB7tqg5AIB2YrG6bkvZk0pLL61ikpkvoxlk
5/QgvU+3rbZy+iYmA/tq2/h62lEZEAwZufGogAx9Cs7AzHiTvG/D6Z8MUdjVO0Lv2nRZP/E4W7V6
rtAsOQ8PU8sMbQzmdwXlz9l5vtrJ2PYgpDYL89vEgXxCl3V9jfESJp6zQCJAdKrgIWkMpOHcsufl
r0OQsIF/7IXf4yasmiDpcMB9fcpldlHCqQTkuO+j11ajLOe1lIg5lutYARxCNNCw8H2LVzznTOxL
QT15AEVm3lhMTgzHU4vcnNf3G4uayBxl5nHWLvUQPgASclR49yQ/68cmuJUXYoHOYwTfveLd4V1C
XyAel35CoktDOA7aGsVoXGOoOa8D4mednq6JRSYhuxTKS9w/1YXGWW8MoTDK3vBRk2LkAXbCCH+h
KFSCdRGqIYN8QdJ0aNbcqbLJ/7M0sC+maXTUrf800N3LNCXc2mGqQv7kAo2Wep7PXuHs+08q2dm2
HW+ifdk50HNrMJscTlRGUJTz4/SJ6ilWvyMk8nj/rF9r8PM9nQeKim9Mg9oAajS+lyTqyjxJswtl
XZs14HgEr9od+MQIrNXnsFESs+J+MfpTVGd9FeZsWE27uX1wr9DC6PLFGd2JpZ3gyRXM7dlTcj4+
qa1SQRDNY/kFHqR9uA61jSXmcqEP5ruPoUJB6ZLb/LV/u3ljWpObTcfF6tq9Bg1kqMoRvaam5itG
g4JNIDPqS/jGTyOTsJT7vyP2SFl7NP+B+e4Kz/5GaJws2RdIKnO1UEbhunq3lfLR4hB3Q1pabUvL
0fD7zT6jvE+oloqREusL9nU8XhrhdXOvfgn0MZgW4okc0qSsVnk8N2QeUBDHWS1Zd4y+ANzg8uVa
0OeqCCBiSQDvYOckAkPna7L5XNkdwfUV7k0svKhXO2e8IhCgwbQhgHm+jyKP7jgJMtjmFSOfBCMu
/A5z8qVrxOleOSk44sfpysWtw48k0V3lMLzSS3zHSvo51TqOABz0DycZuN2ztCtAvmCsnFemYH9Y
pCLIYOfugJLiUt8TsZ/1j/L1yx+RVHb86tM1c6/RANsQLGghlAKX+VaT+MYOZoPNI60ApW8+94yM
glKG9zQkd2YJBtGCo25Ps4eGXQ8ey4UkLNAj7IuGygtgthl3KRHFzpFS1THUzYNC6AW3xrZ6HCKQ
GkGwta+1qx01nnJ1IoTiPV/xsIiLcuvWoIBorfUmhlrbhkNTSCr5kL5462AkuQX9xrwy2tz8ouMS
SUbiRVu6dhm9NnYYlPadxj9XeF0uGpk7J8Cc8ehcewc2qFrt/SzT6zzVZb0Z00qtElcxpvJz78lI
wJthttAH9SiFu6Gt+gPIj4D8G/6wUyzWCop54kZb3mjyQBfZ5GO5t9Etvqb8MMdh7zAizCrUZelc
JktQQbo1OprtIriP8IbsexkkB1F3H088aJycPoU2bePgmsdSm4MHLYzKcaxhGnAul4I1Z8tGd4ms
6e2zQAPYI62QAx5bOqkLf8/oWNnVunIHUg3eiPLTL9ldFq1GeTwmoDsPtd/IH7Ei7UMghDdAqxYi
qJF4f0SJ8tPI1ZsE+E9uCoVZSUSjH7QCBfDvc1h9qsyAjWxo8xs0kY4OeB0DY+wtSJ7B29v6jEkS
P4u5MR7gbMcyTE3YPfluvnFd7NRkZ7r2AAlA9n7JF7+zD2AyBc2Xf7syemXYoY9JfxdgVYR07YDo
igK2A50P+ukBbdRrEihFwZxgJHXp1BHgeO3mWY+yYHJYb9BicH/9CrNM5h9t3O3H5W82Z54rRKsZ
oL0hAteTElNJrRNPyfx8g/0PzdYpZurQnDUSt0rXw8EvkiBNJX+jqRuZ79Yx7nOBTN2/7rE/d3Uz
U6GE5iZ4Dqc8ePjVQ8pRru9NkBSAQjyzh0owlmtF0sc4c51aFsJX3trfKLkGakEgsk5jpizDaouE
Dr+U21a4Ogwn6IQJj5h7t3nyNeY5eCtmH5yv5mPpHp+f493s3WqrwjtPX56CiGKtFmUOebpKd0sV
fkT3HFNC4F34vfJPP8GcjU1e+4xNkbCPuoLVHH61I6k3j2h7HNZb3h+g8J6QD4IKvCvabzmL49hK
qRB45NcvjGgBIVMfkwl5DYeOUtWhqrgI8smC9VfAfhcsQiWoSRp5EDRSH0A1L/rvBwD1g3DdLpzK
sjD+GrniZqKwBnm0NreJ7zXXw2HXSBnn1YKd/0Q8u66gfx9kUnq6NmkPNHaKYxVRLLmV+XGUPZnD
nRk8z7hERqcSM32aRQ5bRgMglEWdpyBowMz2s3ZHKsSa5PCpIqlIc0QSERdZ41sMy51E/tgLwwUv
epXwe/V+J+cRGdO3NMjAZ1dhnSj/DchAWENqLixcj5wRCNkO9XciypdevsNEGlhXqB0NoGWvyuEz
ir+PyuxwbgH4CNLVJAVNI9gwMkNTba2a82taRF08dB0D78b/PN9KkXbGS6IFrqRIO4LxPCr1aAwP
z49UfvzlSqsiZpKWvaPWjCSNyvBXI2Ae/nxsV2RlAIEDvOTtDU7nRp6VXJht0f143NmjWBZQPOsJ
BMHP7lNK7OqQTQHi2QJGOjPm1jcvqP84N0HkwJc0ytFKIUKK/wRMD6YC4AlJtwJmzqCQSn/0jPwd
qWkpPASkpfI29rK39QCN3A05ZeSIQIqgU6Ankeel26n3lVNbZnK7sy1L37exlLeGbSa0++/UbqIU
GFBz3Fuu2IP/WtBE/X/Cfpfr3GJA5x7tuL+xu27d2CkQhu16wTcw8jSX8knt3XgQxGYRn16Cqc8+
lVzssrsqkkxc59ZKsXcmWBdzNG8K/Ju1Bcpf27mQGEEqb4Jg+55Kz9KY8HUgzHQTyrIxdMKRCCGB
UF039ZbuGvhVl8sLK1I0k9kpRkmszf5htLe47ofrVjOQPjYTgjNzW0AhgSG8vq71UrBZ32sMl+sq
Cp0mqbDnTNOvwksp1EfWXlYQbjVpIr7PVsIsWazePcx6sIUBNksF+pvaqgwfzUkQfIvitrWx7aIY
1jGnbYs5Sb3hIBD28/yxK2hku4D5gFfd1JGT3PK+/g3sTN4DYfS+IChREGng6uXK+tf+/2x71+WC
m9gMv595YQUTyTtB41U8DNIjM96bxNtpee9QH9SYRkepVwVDxUJFVk/SAOFukn6mChusA0Jw61r0
AyVqMpSucV+A0J0pPgtFWakDxMV1B239yyR+Wq4UKH6VC5VZl942OCsYCE1faFxjPf9+G+3SBB5N
7f8M+XPtC/Vjcz23tYFldED9d4Ji5o4Hl3YyV9/ZEbJkqCXh6ts4mRMJnNAzojMqjWY1wzxy8fnH
icDNlFQFYwxFbLegV9/46h7XLelNGqOn/bl84NtNhy6PmAma7+5Y9C6FYnZOeAiemsTOzJMCpWsl
qIYltnV872e+RHSKtXR5JZGz3hM1+3gVN+ZiesK7Wa9jcnqzkDbQu2S8EV2wG/NzQYiupEXGIzHE
Fl7aWO0aYQxWGlDEE21lB8BmcIEoVOVxIg5qqTzWM/Toh+lHGMeZzScE4XRxS7ASIRyqk5t5By0R
fQh+RzRpi3LWtMAzTSjJAePD8LZw/T/Lexm5iYdA3rEEuTVh6g6wk/tqaN2Bv06jlXaobA6ky54X
DlIjAYBtlDNOxwUJtjcUD2gX4VTuiFhhVgjkVIpH2jCH2kyv3mD49JhcI/AXmaHtd0uc1jj4ndLy
ZPN5UtX/pFMjpCiMzQM79pBJUTVNkAM4KYCcUiX3KBO0+e1anx9QIl4Zzrn8L5TSzpqEtZ8Lqkag
LmzL3uqY9LtvXZaNQuIlUxlVW/bb4P64SuMMVkUJrHityV/9Cc3zbupDPd4m91wUq1mOwyULhT1D
Ee05F2FOT51+IFPC6nHJYzhGIQwSHaY1LsSmkK0ISH8lkeb6MK+5yHOUVu0vdvvDOITm9PsozUG8
QAbyE5vKlSz/VCRIOSZFfDWDPqIfqEuaCdFMLnh5Tf0lOJIGhQKObWT+VEJs2lfuBVu4Ld/omfr3
pRpqlyR9xjbaxPyvBdnvg9Uv7Jmxmcuxa6CimAwlRhhwcck6HR73OQYxV/ViBr07/Q/qzgILUJxO
4IAwjtxfLaeFuvnfdGWqaYrjQylhKytM1nRDQm9FI9VHh8Q9e+JS3s5T67plR/6Lc33Fi5Lxxu3V
mF/md685/dmY7Xc4jEKvBMMDMRcQNZ3PjknAzfMMaHX2xUPvbzfx6Lr0H7BMF1BEw9ChSeNlbzzr
GWNivfm4xt5/sQ/qqX2Bs0P8bXGGKW/KvRgmWYlmpRQ9mzcLeLZT85IGjDdGPUSa+ERtVcufrHaq
Pi9g6gw4LaV9UAkbd2GhQ397ASBC/B88KUoPTxa7bKshqVuQqMI0jeulMOUMKksjpeE7BLSLfs4d
NhLr39fchHYTayVc8sarK7u2I6S1OmZz8X0076GdvaTalLiHG+c6Uy9+Z1hP7EtfHmSiyPczebrd
XLbooRRE2ERz2+I5sprxiXP1fh+vjsqqYKQFmXZuuxdVM/BIeH6CLIxIgPmLQ+dixW+6Y50RM1D4
Y4E9WmntNd30BjQx+urUcfCPN68JdtBeiMYvcsl1F4XTdGcijZEPEkGg5QBqcqv11lKi4qinN4XI
qOPTzAdvjWpG2gsulxVxUiszgRbqEBpp+QyhkFenHZcC9e0oRG4kUBJTG4T4v5oH3JhCp0DAyqNI
ljjGi2YVxv9naUoZUypqUvELq80dKQuejW/KsNLAQpZwWwDR5dRzuE8O+R+3sr//uSNZ0AECGQ1B
oPlvqldWJYpySJMu4DMEfTHVn3XD2QuctT4PfVNUhOxIiPvkJKyZ69kX+JXrxduvwjEdPDBxr9MI
SYj53gjft857BDDSmPA1aBpZk2bCC3RSvmA3ThSHeHn/TZeg8GOw2ie8XnELgnVDKPyEmbNd6vPo
j03hnCpZkIvIQyXsIRWDdnKeJ0xtxWeJtb/ZIl0bvYxZRNAdY0ibvVfMqRFu8RQL9M4PSbxiFnPX
NdgFtKzRVmwupyy72AwC8ZrSX3R7BtmTyfwFm6hA/r6NKXlzcM1fknKa4JpsGwJRZRRjPgsOq3FK
EDv/z+W/EIF39q7CIVe3fL2Xa9x5CVUIgqicdxyqfyje+LNoV8K5hcKs/qC7KkhgCxGVH5dDHKAu
fJpwaYl/T51JY8JxVNsmNbnTjKud01imlJyn76DebI73JgWVkuyJoBvSl0ltn6ypZlTYfdUfCVdR
gNoA+A4ZOkxQ33I8DLw65p7rHMsbJHBdttQgg55EHpC6z7LKRsiDw0exvNJIDeqXsoF7Xe51rcYK
Y+WA5C5/gOSttg5AAKNnv8IazgtrAMbvwezJ0e/UipbWcJNJkDqY1wEhb3bfE8TTi4ytx0//fjQ5
nbb0/SoQIJapIp+hZaGJgwsCwaLfmbGxyZ/UMrBAPU2ir5mDJQonPChdTkyZMgboACYm96XDGTRH
Nv5q5WNgyDUaH7PvMEAReJlRpDIzgnqxV4p9er7Ah0lIb78b15LUTTMnYj+wWLWOzKzObZ1D07vP
5iexQ5XAvpN5Kff8qQoilYArIax8zZx79c/d1pUc4g9BDi29hdYEg9RI04nlqW1Djfq/lN/Dzmmb
V9T7mAQmkmbGxIQyAemJOIr/fWTU+oYRPaW6Up3AlKt1nyKCR93MJwU8C9q8jYMiUPF92YBC1VDe
7TOM/B++5+jOBxDZqTm/7MzplT1Aed6yAop2I56LlUx0FZfGj3+ecIO39MvrvJz0zlN1Il9WjiKG
rvQaJyrlGT6KiP+B3ApLMXZa55w+3vsot/sBlIzs2waTaxMN0oskYuMoYG/LngYu//v/5MODAJzt
dB6ESFWafs/eJtbJZtZ658U1qe2s99dezGBpccBAQ/xc8t9NdV1AE2B3ziTaqHOIenqhU+F/HY5x
+wiDNEi7SD0NWA/YBFDQQcge9PH3UyUTa1KV1lLEgvknDdizAsmaitWsuvbw3Az0gpDOmEq962mN
KCcAWWrc+bm6ZCjnE7YOQ2V7RNSd7ZauS/CI1ycy853MMJD6wFajHiajkFcHjObw8ZDdXzsWaO/m
zeBdoDidaZzSwVa6rayp3JPgygluFF0NDstBcENacUk3XmpLUStn9qH17CM/2GwMd9QXRFXre9cz
mpvIGAVqA4+u+zr41SpoX5WGkQGfEjClXG7vSGSVDdb8eCmA7FWs61lCS8GvD6U/BV/h0sExfCWB
FS8jst29vMrvWIBSl4C4QM7E9wtKDcOK2cS1p/q3jwQV1AH7nJHroOxAc5lh52Pd7H2RqJezeHL/
wJQgVoAe5KnyVo4zwoYJshXcDH2tpXkNVOyyElAWDLvzlZacnjWPTpQ0PCIm5WZt6GMDGh1MXm74
eQhrsdVP+U7UWmGJGLJu+DKmlXJ+7lkflJxJT/W1uepMmESE5KiLErLRGp9xkxjp8D7zouN3QGzY
JilBBCN5bZbpkauvBJy4Hmhii+C80+uCvhufn0Wg5zEW5KvKz6XkB4Jr1AKKCwomKQqz5/AhZSrf
TAbzmCOR86gLQw1FcaRigUrSGWOEzw8q6lAhOupWoqkNJmFYhXdQAaVLnR1XubtAdl7ieMcRKCrg
No3O4nE2caKV+b5QZnI8D19iBeUKLVcjTTqhUleX2qjXAjPA+Vyb4viOJ3sZMOYAlnxYno5ZQHuL
FlCZebWoRI0E6FzA8mQZXFNe+6y54rEv4p9x0jYG5Gz+HFXS/JUjh4i+4SmyCHCHgMI77XXacuwl
ctDhSpwCUtRs/WFurJ8V89DC+XZS0PhhDjb+vHkKZzijqxJlgBozTJiiGtX/9mmPfoPUALPXaqc0
HLSuw+ahpkC7WeaAkhCpL7F+6ToHUcAtGclQNR20/CDWbYFuWVFnqF4mLYH8dgmjDv7+Qg5L6jn8
nEt/RSWYaKAl/pXmHUxvEcV8WyihuUQUiPyMKRquZ4p2ttM6xE3/hzkpq6XMr25ghPWhXGpaCKWv
lmLwJfmY/yV4tLTG4SDHoiU6E3kO/MnqpAQt6QnvnIPqUh6iobKiMGgy8qL3KKioK8QALaPqcODs
5BG9mZljKVSDy+rgr/UpdvCKpSEMye9v3x9/UFMgN1bNLHAcYMPthlG3cBTyKGK/Hy3fUrJZQrmw
KWGrJRVda570hx5rvBJjM21drBrSa/SYvz1+Ny5Z+H++yWGv/6cHtpE7Bg7GyEa9+2QPv39/DULA
cxFdRbXWaxclF8GrlH2bTGu0jxjSIaAfy9nZElvVvea+4aUpNzicad2B6QpaMvpcL80Vnmidr3sY
Oh3dY0SK5H93VMWehSYZ5JOk/4Uw1uU1q0+fgOE8SlihdCzM4yjCWY0gIG9tNkJ9yJ21EHo6Itj4
CwchTOxRgh1sZ9YPVH9bs5ON9F2SvwH3bcVSCYsVs8ij72BHZPDrNNuoHhjLKFzIZlgBrY/ylwCQ
MW5B0PsFET+q7gvJ2enIkwyThsZCLnN2OAx1byqXNvVg+2uxswDnk1w1uFvJHysbPcMH5YvPNgnB
RNvMIsz7OEkZM06OT3b5DZ6KpBMz6lpSn9xsEpD0quwg0eMm0r/ai1z5M9bBphlXpcMwBCpoigfM
8BI27bdlhwlT0C6/lGXuPxNA6cBAKCNUpu/TOmJbVMD48jt1Xs/taMHRL8mpDMQRq4p7TSvaSABv
B04QREuTd0M9S9/3hkh6XJmD18AWcMNUr1Cs0NnIK1qLkWGfrPq4prAzfp7uQohhR2l3LCyhhn4D
PZiSQEZvxKgx8r+lrlCyu3WB231TupAzcjDRbop4RxfMlxejqqHvlVCs7S90qLW34D5WRcKDPRTU
eypbrfmA0oyboH7MAAK2uSoB2/X3I6KFLAdG/L+VSY1Tff/2enhOixh8jiM7Wh8Iyi2cl00P/rph
rJfLMBxa408lEm2Yk3HUZIIhsoJBJzIluokqOQ7jDl9wxZCXhbtsDgO0JHbIlD7UtnHnPhjeVIOX
witvsFzW/ODIVZ+GIOBjL4eBv5fqxMQRQ4PIvNFoRcS1hKYkSwVjVoxfBEjU7c5uJo/HEyGV6P4o
Pe8kF5jAzysL4P8EsZYubhGBjNfJNVgDS78mt0yI2GTcY016WAWGF2LLzW6gpx8nU8SSLS6r+iPH
36+6FAkvnv1dRuFRWAvi2P1Ba0NrZCpuBFC8rwDSroh+O7TO3/2CQOr5vPKU2Fi6Kuqsi9XGOc1g
BBlD9jn3GEczfpowQbTKKk3rwUFQbULbvlCVIbvyO4fcApydKcB/MpnoPkMRGRwIrIEgf1fA380K
thBsLPABLQjDHAMUQo4Aycrfq2Az9NnH1wFsttBk+zSJW16V4X+szI4egg7Lg5PubOP6m4ZB09La
Qbeo9QTOKeTS7hvGyndeM9qBk6XGl/XMGoqkVEyM6tkhy3enquHKIonNMFxO/gEGwRZaO7V9Ip/i
V373ECFtqBNrb3HX+EcmhgJbe2cBAKxpve2ura0cL0p5/NwaUZJw8OMINEaPeTkZnfrsq/wwv9k7
lEM2WZOfdQzPSYe04727/tJyfF6NFn+yXHPvMWzr+VARuPmGB6Umh66yrNvaSdU6KSmMtX99QaGj
FbPdanaAcB0pM34E1R4yUK8Q+ojpDQ4DnRJ7KUe6ZzLoO+yHBl71wHyTbRrEn3g6ekVh8CcZWdqi
FuKWQSwhF/WXmveOFNGocPkppNFmS6IuPhO/li2W/gwe3X4iCcyfztXYW5tasfPUk+vtlWmO2Cxc
bRViStAtqzkPyaOP9Fj53uq5LdZTSiVbJS+zfy7i1wly2BJDCEd/PgPOUNc6BPfgFpAqhI0dqvt6
dEKxEUhnSqkO9P5GMl9SsYUinRi1hyps7n4XlqJxAxGKVnfNtp9/hXaneE4JK0kRJHDtIy5OtK7l
XbmOoTGFdtlOG230wLorHdBfWNXasTg9owoNEg2/kzgiwp+8V7byYBw56OoqfgW/b8m4QZAftlml
wPFcVcec1AQNiqdhM3N81mqCeM9yfJTXTHe8HaNr+I8YroePzjgy1l/lUnO2hHBR0Vrs2GYE9Siz
nTHxOfyaUJPxB8gpKZnUj0Xrb6/f17ssrIWgb6JVoYTUYbHUGeQSJULGkY5NSLPQZbXAG/grt+/0
zrFzffxrSxgv4qP0Gc1KnCV6PQn3qAJkJbufcXyJ7SGopi+lzJEc6xjyjFSGNSl9PwVClIccCq4t
FbIqKMPvajI6s4GiDUpzHk4XHAcq5Sa5htN1Retj5Hwcaf+C0v+/LH4dJ7NiJTCNuG00C0iBw4/E
ouUDMgcm4bfgiaI+PUvkJbkwJXbDnp91FvadQjf2/1fznlHWuOfAV4AW9Z1TD/fV6SGz1JtTtrS+
jUbkZI6pkH+ZnA8+lHT3rtocUxAyRE1c232Bax3LkK8SgYyVD8qQGZvgo4HnDn1aP0DdypjjgLHg
gx2hBuAxTC/eh5YU3wgs2yYT9ZSgQipn6pNgv/h4xGxAXeMhlwRG/JncJXYtuewDb3TDZq7kZuHI
026KZlPcATVE7WaN47rZLYmgaO9qjQ07KtsVx2hTtg4ESmQfAbrffy4X5vQ+rPH8U3x/JxT7OP0N
jLqVWZr1BskRueQExIq3jLPvrrHu5CbNZ7UFk9+RcOMqJAmMHM4ZmIE9R+9x3GBXW2cQPOU8OYoL
VOHMgFvTGAkDw8qSIL9r2iyDgsPLwvQLgbKiFCSPv/SP/g7tEx/DbdOPigvZeGCpJsD6uyV2iAuy
m+MBy0ds8IQaJcL5u0Y567j6Dnp11+MxQsk9DBA9nH0ceL8ZMjycBpM4DgenAzRP78FNfW0z/WwA
Btftc3p7vgJfqLC1mtplrg1l2bumN7poG9CuaySwf9DlnsDAE7qBLEJM/gLDg04i9TrfkrYRts9x
0Im2szBHrviAvZHDMlG3s28UJ4fQ3o6j51hIyty98gPmD1RmJ7FKvwK53DoqNUFvp5Gvf+A06dY5
gJOitkQpe2WarJtli/mkWJWf9eM63q+Mw4qbjNIyV9z0rF2u8KLhuqEgbnWOHl3/64ggyJOz+r2l
odXZdsmCxnsNUDH/AzGKK1PONGW0p02LdqYlYzW0QB0eyo4OTHHRYrZJk4rJEm7XTh2nOv5cHKqi
n8ODqngt8uf8M0zD01gZgv4k36rCGIy1s3SZ9PaO7RFdebTYf4flXRR6IEx8R+Ot5356Wb+hepgp
R+c3OLv5xkXLFzt3ygKRz9wyRNYWv4AmttHM8CjcChcs4v+YKkqa8B+FaDNm+zh1GjebaRguijwM
/QA6qxV+04I4m1XJleBddX5ZWQ6v0bXNAU13gd/f5yT8foqDgfJGW92Jgqve+aeCXcA5gbu+lZwR
04TTrMkUsVhKUTNzl0oftx4Rx+T4s/sjI9GZLZG/WJLgnzt30IqgIvvNbSmCogeZ7UmjMpZDucYc
spK+IV7H5yj55NILu4S1HPW76tciLIG7PHD5xYN0xDGFENCObjAvJ+VJyNNzLW7sU2PbYt7i208/
djbitsiNd7Ld58zhelv3iOMWcH3QksWl7w7rfcuaDOoeCPUU/2KLT+3Zq83BmJHWJCalEST6NdE4
z9Gt2v9YZOaOp6jm/ppoxc/gXYubMTnk87PjKzvCcBY0kgEMMrsyy9wdMTxi19BBO9Qe1QeNmIOP
ftNDCneSh++fcej2X1diD4SVpzbDbLtSaEXI1qiOa4s80B3bHVN1hxoPTD5gyaSrrJVMaMkgU+9T
wHAfblGwvSc979spDGIX6XxeCQgPwVdHjyoYAZe6GStfiR6Zo62vd53W1LGsHj8brdaH/EI8p+3e
Cx+bpXfxWk/wtvRWis0m6moboDf+xf0xeoMmPcqlOMTOc2xLsPcUsyEJz3xuIYpShsHxjqJpWmyT
kWvoGq52mapcUD5Cd9uCW6Ka8PNzy6zCVoMZSiGjDBSxJG7Ckk3VlR/4+BSXERsZFEPibRBc/Qmr
HKuhkzVrvEfU1nwoqDo//lq/F9Z/+FruuhE6pOHoggxVdvnbjgP5ppsgsZ3BcpbYmCwckhPfWmPB
7wbWGnBkfh/JhBtBx8pDV7ZddKSUQ8EwMiLpfHEWTgKwvvNJqZnnzzlEZFNQi8b5FomUpbefs8+G
P+b5lzkoRCGxLP+gs79akY2I/4v2PlL32ii1fSOB7Jrdpbs+yq5psPoBwkmTZT0ga00QrGgN4IDR
xeb5reaHUT9TZk7YcJDRBGRMpZYMWxPHaMpF1NHfqgntB7nng0K/EkOU3EbAppja4+RwTDciSCll
i18mvz1FKxRwR2XoBVkQwq4wjBbQGrLKgMUVgBsevdcLquUTFAez/yck26lrBDzj8/VEnSReon3H
WJqKNR88BleqrGf7ZGHDjKhy4N5zbF52CqWBC+zX/R97A24sFlNWcv5Qqgi3bwS6Qf+od+VeKcND
4pOIDYUoOuMFd2XnzrWm6Srz8L0YF3jV3OwLqTnLj9eJ7OT28Wy0kFdoZbVQ9SSO8Mhjf0icvCIK
xCWNT41NXELR13rKyp9Yj2VwNpB6KkeN6f4Hwq5GkaDk2Gsjk5gksOSYjlNas9Q+TFdC4FPRNBk9
goAvxS8jGHUKyGm9v3HsemIFGdfvY+po5b4P2IsfdhpB4HO3KCFyYeHrpIW7DAgPRsFEHWQdkMH+
508EA+zM6TKKYm9iN/qEL1KoX6r1oXZ09cV87MEDlKz52cJHD9UNVyNAufmEGzlLsopRS67sHBNC
VVpkU8plbAXCZbM4Tzy67KgS6opvFf8UihTbTZozBNzIpzQOqzC8gXuS/U1T49zcqybsOb/rpQDS
QpM58aaC6t8cwLvEwmfEoHcTQ/mrWHyKSqkpZbcX8CDRa5NxCA8aqs9CJCloa9XGHeffDsNwstCa
pt53Kcz9FDTHec7a7WEXwUJExV6AjTMqsj2UjYtptx4nOV7lZEPLKzJaUrzCyNWghMxGwynshgwo
aWtYVPhtA8sH33zr6QtYgzNB+wasC/4gzKu41lWZH81lOLAaNoxVHd0u0oGCg2ivZBgNEAtVIcsb
im7n4QOYaPvrShX+0I9MZFRG6VHwj+xvCh4MhUgrtxk1UD6T5fn2OSMViSOkZsrNdjO/K6ohsB+1
7ktrYh5EHgKuWY7oBAKjfxUxAt8nIHulqSpat7Hvc0CphlHzboK+LJazAEM6+3LJuHVS0T6hOMGP
mx3WFdN8xRaotz0XeUmH10vp2fW6NxD2SzBeDAvfyQbC41g82+fpfH+M+0h7oORz6yEi65Lb++Jl
F5TeLz6Q/LfzheEADxMnObWUg5dwFkX6OuktV4ndumbzZugPKIbfztdRaxWktycCu9zEen1dzohx
BFZdLAjARWTNfa00+iHscxZcrqknt47EZ2b7IQaV0tFQH+tiGKAAVuUMxcBWlDpWm76f0GLQ4jqJ
B80jqhZPAQTZCkzMh0EYaoC//n7E9Ed1dZZGEbV1rAZ6gmAsihscKVhQmQ3t5r2qkfoFTtqRbpAi
p0q5CDuMGiKMh+ehlEYHopLdNYieboGHD0KeDZtPXHwDDiwsNIQi4QBL/vps/V7uOgAr4q9cn7s3
U7FogHafHT1p2OBQjnmvwIV3ij12vLfJad0mta4lFSR2rivjAIIEd4Qm5C++6stXttGJK6nlXBd2
3U5dZf4/1txj8+PcuGeE53uSX1l/vrFhy3oZ67h1TXPe2d1mXmfBhspidT52rBcWp62Cf1a3er+j
L27h7te5olyNEiE+om5a9MRPae1fkTI8yVBdjv09J49cVUqVB4d7+AnAf9OR19rKHgl1AwR5vpF4
7kX6M+/BoT7S8LNfmwUBe8MatkgIcF6KgbVWq45kdehSuJ193FK46tnr3H/LBP7T0J8iTUmVZ2yd
e9G09LjtFaLFUrICemcCbFm08KMI/CMvlHOHCWklI/ErrsWxpuTYEVfP4cnYpiYdzL82Hp4lKLfX
J0fUBlMv5cx1Er+HGPg+9mM+d9Hym76bpDEghJm1yH4xJPLpSX9ynqK7wOvrkQ64I//xXV+OYCba
gbcqQ+JZSxSZdFJ47ubBlJcYwHqnBTWazxpxnNx8yFoMKBQ9t8jK4VNWp8kjMyOxEvJOCLHsTCOO
cJboPmx0DLjy1zXn7A2DcnoEUJIxKxf0LxqpxuA9R/DncwzRXbrkIPw2Yp8gxN0Myq3MT/+TydT1
oP9JjE57GIg10dJi7pIZ843kvXkaO9Qdpbsg3MXhcUzDFBlZOKW31Enh3EEhiECNvDducE0855rG
A6xnCgZsDcMsMWecv+v3oA+eT+AdJKqrQf1D1XDNDvUuS2/30qCtK3Mwl3AAjE7PRBpSpo2B4nvs
ATg8fBL2qy2/NxH4Lfdb7vWYD0Y3I17YNEc12IYOqv0MpHNXF2F+DxVM8RlV45BmGsgQ3i3hU3mI
LYcFx0CJEy0qFZgUkH0k+X0hlYbPC/S46is9MJynCwjdNPWu7BzEDvkYz5mc/y/N3+IbVRrTXM+l
JQznHmzmBK4iQEwQ3jfnlMSwh+qdWSwYdSiOlzuKnJHHJ/+dTTX96BQ3eKiXOtrCT8Mk8cuH1Flz
XrxJ0I8pZSrGCka3Q3AQ5H0qjsoN8siB1nUNoAGWiGKLKP/3jUAsZPOn2MCN+iC/kUuTojeM/Zgi
1tx8hjGcE+Es+vwxIJB93jYaiyhxNjamxl4cT+TGRW+4jGOdgpapAtqn4L0xF+W1HXfrXf/I50cL
8jDviHE9dWiYO1uHaHpjCnZWmNCOYcLQcoKF2mVa00coZF2d77IlkgjVip9XRgdMf6F5ISG0EF3t
fy5744xgjL7maNVNpmq8J5yX+8VYoPXLsRqsSffiEONldmML1mWiryzQuYfGui+/hYvqi/zzTYaK
PYQ0CXApKPNEKBt3YZGOgfg51AFG/yGWpbNI/hl4BF7jJxjTg/gmPF4QwmsfOODLaqBnsbYMSAAK
G4aGdKECpAJ+8CYCxVLRMZ/62/dUQ2oMqb/9jUlIdTVYm+qdAXLz0bo7F7Zmb0L9UrmGetM8n5W6
68OPv/jQ7LMlDQ0ZuE6tz21Tn463axQQTGbvJnv8G0WEm+mhOtRd0P6Nd4gsLpiK21GaRjgHAXdX
uf6rCg/MG/2kQ653GBd1eo/jHRhNr6Ysro9VRXMsvzzoy1pB9XADw6sjJWCoFIFIE8DoN1l2+JjR
uYLYskwRvEq2DoGszSVRsz8DkK2r5Mxwx3GsgxTOQtftMIBX8FAp5BToYC19XjYThnhElc+JZf2h
ViWbq4G/HS5kaXsTNF2lz0pBdf2+ceUnMruPvid5z2s/HQkwAcL54KqLp5iVqt17tsyH8SNlJZUl
LmNQ+ypBmeTBHPHqNpRov1SPTAmx0A40yEDyYQWnDPyJkNhgpFu1tqnq65E5kHpkXQkUr5zcnzmd
teMcao47axwvxK9y4eGgNieq9UYZ6cqKoeVQdTiuI6PJMrgMdJnVFwebBoRxw8a0YmooOA918UrR
zqjWPcP6H9HNMVVRnMn+G4pZWV2oUvLQ/lgTfnWyfJ8A+qgG3hZ7p79+CBNuG1gQKbHuH9MD8ZK6
Bc+5JsjkQNhUT9vuPGRLc6Cce6a7ygeol0YBHHpgJO5yzc99mFkiUmMuWibt4ZTy6cgxxgwxb5by
Nq+MRCgM/hdrG8y8DnpqOe9Av5LnFwHiw8W0Vy03uaSx/GxrcOuajpbuRvt7pyjYX3il6yiRqxch
YIkYb2b7sl2hBEWVBYB80gMvFaCbVeOlIjx7ZoYjQRcoLTN6jFitIEi6uLySaWTrveeOO4XFkHhP
qOHymu+rYT4aIZYJq3+HVIqxDjUbW/Vky2I8PTQFAMpLPoYosNmQqMFAqzco4TrFs9m26qjqlP+V
TW0OosULuYS/WyfvECXbWc8LD8+s85TF9nchbmTdcYheQ85d9bvMp1Dgv4SKyQUu3YBUcc3Ye5wI
9NXDOV/U7ieCUyC/4TYgj1W/LmIPoUhFvLGqDAAnzs64q1t8yt4G/DVzqW6SlbixypcOICDKR69B
F7+4RlSq7iaD1X2z6i1EihreEIMES4tOd3rlQipTNv2xAoJ1A5xhWv3E48KK9TWuqmPNXjEQFQYA
CWB+mLIq+EdnvLYNlASWYbTnaUea483XQPAQtV4/537TU6QwAKqJH29AQqmhdeHycloxGDa1vWK4
Io3NH6HaOMd16HNjpe9l0++f2sk7Unj695aKaF6yk+wly1H0Uah7FZcKR4K2Z3sN3vP4iKuGcvfH
vOGqVrOmq702+eDDEBDQfQ0Pk6rXd7HjqQlNQGX0vKP5mmbyqyuVZ76wvDn/KSKzeopWz3H6H9Eo
1C1cpx0B3JBhYXXHp3N3LbT7ir3lc013t/RSj80Dk7fljMyD5UsWvPJhjz3tH4mccQ+HXdLCyGu+
rnlRTlF7/3G/OqkjE/uarDUFIYNjEwAXpTYbWG094SHvF8IVzBIuGx5k0+SEmfzPyFRWOdL9IYyT
nPqAa0fJXACxPdzzUJvv3Py03l6aYSpb7qXr9y/aCnQuDopEn2PFwrILDJECJjj+9LoJBaRQrX6b
CX8f0G1oI9Olxlhf1hZlz0o3VjCefRRG4tP4wE2889RzuziuDoCB4E01K95VUH+uaJj77Vfijqdv
54Pi7id0UdpRQVOIRoaqXXm4+vyHUmBu518iR5ZyLBKgSTOks6DbARD99ChC6SPXuari0ccQWlEo
gUqlKX/LlUz5p9xhv8A6ggpBhFNxC5DXb4nzzxFYDZjN7V7XnICBchWdkASomHQDn7OJ7/zXttS6
zxqfmS0gh0s9CLz5AzTdnLzcFF4BNQlKBE9XWADwSr6vqNPwfT4PEMSqkmTeKAop83yvZzijFjyx
t6EhEf9g7eUHmt+vTebBwlBrudlOHcTpocWjwiY6GCONW6I26Hegg+6AfZXBf6TvdohHfAqqNk9Q
ul48ejcDX6mM6tO7ZEzhSMHQjWf/SD8c7beFgiEQbBNP4V02g1g4+GHA8rhLeDgctdRQ3wHypHdl
FxuhxksmVth1JZrEkwR+tjFLNGrHDMxt8kQ8u49MN+iIatPf1BPZ53807NCwcHpQUb8pk/gFXMxo
n5c9Hj7KjVtEgyOPhEEEIYnapP97VgQvGG9HiASPhKWtSyDulzJPKXx+isAlP8H/r3HzNgxuKoDB
abobWVtmhnoOfew0Q/E/smtkN8m2nUFnvjOY56jSKo7ggvmju3TGz0bsU1dDe9Ktfr6NAP9ICXNj
BNeZznrYupO3Pr2omDFT0Ga1joiN3nrLm8PY++16+PWItwXv5iHe31bdtJfIZf4dpWiZOHiBrBcR
agT/AUGQRmtqWb1uzp7t7spz1xGenhSgK18neoRobpOChdPKt7dBfxZBzSiiQUbwr2gprD0RAD8V
iZ+C3VZlP5cWdnSOG0qbWtad+gsU8Vj4EXRJv7ieAVmAyFSZwr7inmyg1OGOMrfwUNxxVkEJE0vs
Tf04hbsx6Aps+AvsbudN5CeMB3A2FeUyOHk1cn7g6dAL8ZuubQG3DSsXe7D/tJ4xRdD1Ho2UKTlF
C/CgfGcaqFvEP//NrKx5paKX8txpntRBTwfuI0KhbWa4GSwonCIfvHocyu/QM6x5EdY8tE98DluI
SvIbA0L0YsPAPiQ8Qn8yfwc1cv40LQ3j1bo7jd4nUswDx5ZPv+XVSrZcQJmmcm6kXoCOTEmtaAHt
8WND8VRz3likk3TVrR3e7fVZsaTlukT0XfEzU7OWSHdre50gWMlZygFd/QAi/sM8JN4vV9LSQJje
5Yb62PXs9/kiywbNQDEJaXHx+aAxrsBEgjqflRwfUvLOvvtYqwuiuoMPc1L5gEG0/gSwWM2Yb0hW
8QRgU3qoQ3dQWoSkc2b5D9vYt4eZdXnssZlOvPAv4LSKLgB+f1FXcJdW/KOH4hCP8/gqAucpc1Na
UGRKg6ceDXaGs14/iMrxWoigiIe18uefRIqwi7unzyQeTZpGfDYR5poAw7rbDVJ6iHG6ifQwnwcg
3tIK5xitr9a6xFawLRuE3M4iMdrFOC3+ONQ2mZbCjZX0CpkekZh8cAfBRn4cWzBcACCz9czr9/g8
S+4KsQCbK36NAMy8NDeSWS20qY8R5q46UA8aLj8uNEIPaKlmlNm8OcEPRwX2E38WOOyrJYf/k+nf
AlwcjNg3o/7A0mI3XAumDNpiwqpA9+Q7190odoVtT1UQGyB2mH2yiQHEZ6Ucc8la5E79dyCfXR8Q
pveJn22dpaoEC//i/YJJoHm3/o80EPFKsg+ZLbH9pohANQY01IpYz1Fu5WWJLSY//RsXnGAt7aKA
/kN3bvlZmH3nUmh0Ah5YpQtDKRX5c7mGGAPj41xaSuSuFLA1I/5heD6z4SMV9jlgOVQ8Ks+to15Y
9qe5jT7KyVp6RG7PEqs8qgT7kwzGrIncPU26gFOUTSE2+9nAC0evpHsQ9qg+c7jR76iCbjgNfDuw
/EYfuYNzSlkzoktJiJdpLBFAV7+OuYAalIikXx5f0MwfVTQkqiYRjVf7fLObZW0P3xjFY8tnLgRg
47cQ6/ny/I6S/HY6piIcGbW3aLHR47XHtP6XVT6suDIxN3C0JtEMXniaPPnAb9qilDBFhpjNVaNq
RBclU9xyl/6e/Fill21B0wHjf4AeScMdQR7NtP6VIysiUDU6Vt8IdSJCIoL7TdYVrytgzQVJeeRt
ZCQy6Rsd49iZ0Ft/7t1tGBEvX0JASkATK8rssZVTWIInH75s4n6rysr5hSOnQywjUP5KNaQbQ+FB
QSl0CjhurIYIiXhy3xwq7ARJlPQRqtQua9dx//DmYfJBotu67svX5BiJItMMBhI1BRHSUbDWYWq7
PDkouJjmEYxtvuMUkmq0o83YH3A5SdUTov3kiVY9WwJ7fukDXMJR27s+NPQb89lFB5wutt9bwZgS
iA8wQ39UHi6R4x7q+dRJ52XYpNcj+c9cjAGzAztaNklLztGNa4tqWMPNhCZKB8zu28p9KDBqnVtp
zqPoSHWecn3XtdS6TN1MPjzf+srl5HlDdOmQMvWX8bsLDec2lQBeqe9KD2aoN1H2NXzD6c7y1hRq
kqVXqfeqWr8oSkLfL6+v82nnIv11iNIv2TzSqTlPRlA9bvwv4H4BX1VqxT2VCtZFRH9wcI7nI/Qo
yU7DVUCdnZga1xArEFtn2LUFbHfcLlsqBm3Cal8gpCA+ID2bcQAbHQrGLQqYIFG3gh0jn5smLSet
OiyHk5sZ50tyk0bSwPKQnePdEKfbZBXXFIIeG4I+rpjIsBCwe/s1QAafKZnjfEsM6XEUNBAtY3Sc
1Yw7pPa1Ym0rCXDYPFF4Ehj+XrPiD7H9ZqsR/4wmCiZgL/BvdwEb2v44kiRY1PSLJe58KJdFV/2t
9WsVeSNuwwk+SIRhCf6TsWB7pYyr2IYz50iFZ3+8g9C4oIGhl0eCBgIlIyRntGDkZbZWZnwZf/g0
YXALRsNtFdRk+FowOUDSfjspg3ckrg141V+KZrzQuqZayT5LCDbpRzvas7kksxmaZhQls20BJOEC
Hn3IaWeB7hHHFuIAF64LIj6Sn+MOFbTkCOKGWRgdUuorU4/+8e4GLzzARhID4FCmP9gvlEtrGpgH
LFOO3k/d/somHZeciuMAsiwNrC+uhdvIGeJmvJ+zXWe7KchWjha84C/55MbaMJaUi671brtslV4a
ifQgKwXSRDc+QuPhEHWI7yT107PbSi0q37CmtNdxrnJIzIjqQfhCPMDtPN8Y53NrR29IhYH5o+ES
fCqLykt4sBDU+WQAkBRgzSf67hYB1LD226IsPi0hz7pe7mrzPSPSYDCFfudyiN/YaG4aUfzeG2dV
CiQLWV5+PQiNrUN20kVMejdWZcChQYBIQhCHOrKJqZPqtoF52Pw3SaWc4YdOTw5tstWPZZeIaoJy
HZuHAcPpPsfW/VG+rTEjZtV/bZQwklbnkCJ7fpz+IxxC8HzFkzlRA9wNmMoVlq4c7tMyK2KdDkPM
aWAY6UqCY7CnCxaEax7oKSEmyBUJxLSN2Fd/0tcQezXTUPRbUGDBGW27dtCBj1P53VvhmEa207tR
AfXDWw68NZZydqzXfnQlkkDGrqBHF5HOgmBHJU5aFqxC/26HsYX/F5PIfOf7w65A3vL5HzV8HXiM
fV4zgFm5Cv/t7ReH5hndwPTQx4qWdjm1THkkQ+PMoxXikGILB2SjDvAbWIkff0XQiNVuSdbu2f8S
Dit0GFapWYywCxKGkuAwSOiDOsREmLiKB+Gw7qxsgag7QtcjlKUEzKACHgMoBqmGJtlgECyNKTu0
wxInCDS4Gz0ki00Rwcd4MVmtdJLpKIwlIwm5NrhZRSTyChA8nGBFIICIHlIaW3lZXmKx9IYNSr6e
7wTE9tEKnCDxAB+OuVK7e2M/1PwD2FYNgo957wrWML+KhHSGp9KL/ChyoqnDxahzIkpD+lg2QWUi
hPJRnljVUMIjkPDOZVKPTGzfOe8xhMfqp8LQ7tYYjOva4otlz1Ov4fbOQuJbN+lwgKE6aYBntqpp
413XsldY5q4lbg7gtl/yw1N+ccRqgs04l6uUZnpNKJYTJNu1cqeXVE1MceQiICjT1INpjbCkNaUg
nDkEnT4Xu3ORvXC8vawY9t+zvhGLiFOb+hfus3W8MJcxrejscaQIF1TIcRrqpNRJQ3Z0KV1mfLDX
CK4hhh1716SQWVBQwVfHX3aQam8N79nW3jwhzrZ1bxTD4xWiuXtr9uIMDCtSDMVxDL2c4G/0luon
uqSKsg8nRXhuyA64ayGuzRLEG2RTGqrRketrannATz3BotpUVLVlHewwn02SXLFLUMynzYAsq95o
HKnh0nQ3Uo1/9cmy+2/NhzlVDebEJDxZ8OfUgNNxfaIid7SJJOnhkc7dxVLC/qTo7XYmdRbQO0xP
0lg4lhRuugVuUfzikDwU/406nYLTWhiTSYn0+l3UJRK3uD0FaosPHyt0fzkc0om0yIMNt/daRd3d
P6ukV00lzucGCFtV24e3aMkhs+nSxt6Go6a7e/j13Avx8liVj7uHsSh2GWBFflxLO+Bq8MKVVYXm
Zs5k/pxLoYZUIdiMVMOssRBT/HPGpSkkugqnUhQY5wKCtiaKn+8HTdBACHVROgPOdgMs2SlLAWmA
xDCccbGw0f3Yaniny8k4ZvZc8RAmFp9s9HKccDsFDEU7saXAh3215GKG/pdc7Hg+l9P+1G6Mneoz
kNVY7pLyEfIXOjD8ATf+wdYmTot4cWI7XEpzcTD0e/j1gk+z2a+xlMf3XY6QkPgQBI3xKLMNKe07
AZSS6M4/jV6iwb2wWKeA2HcQtgarzYnL6QwpB1yik5zvQGEkMOaLsGQN/XbYZG2f9ZiaZE/KR5Ya
ZNf5cBcKTmUsA82aJMQZz3xPGrP2lUGlA9zonSSAT7+bmIN++uLYo/p+fXJYqaT1Ix/C9r7qpd/x
pDjVJYtytZH4x8hYWeP4aC/9YeAQziufJu1lsePesMfn7X8h8wRafhutIcYfn/ntY9kmBAYF8Axp
wUMCvu86quxA4HKN3j5giSPIguZkCPPLsu5TgmlDjGMGusTUYAxoE6j8kqSxLWzk8Ml4uOLhsni8
blXvt/B+eklmnNsDmxfpy7uXUyJopHfu4O5AB3vT90YsxFc8BCtX5JR7kH/mVaZPXfr+PrW2dxsD
TfXdAoMpZKzwSDIkdHwKJgS+lEelMxIuz1yFEZG+TN427nK3AObWqdrQNYrOxdOPhmuCB6glS/YD
V70rp4UVQIKXtAzwv4hhAA1KQyneTxc12K3hf9Dxp27+qbghENJD5GlvjdOYn2lZ7sE0g7a6cUSc
20t4MsbPRaEsJ1pkjESIs39Et5/SOXUiWRUJ8id23nh5kpa4IxDFOQNIXEf8Fi9AacaxKFX0mUik
l6kIgdiOMl3KGs1rPeysK7nysuQvGj+hzNCdFI0ePBnUtKrzBSO5jzCJReFKVjDoqj94EPSuIWl4
cHDeZInJ2f0oCWxn7derAzMbg7mhZR/5D3TBImKiKMsFmEYBgwXYkpMEweeHWMsnacAdXyvV7gEw
BbaVj7TA5vKqk8LfUlDas7+A0HT/PTulaok+0s8yG2ZetqxFrIqMRmIIlns3Bqss2+XITKEgDR1F
0/UW8mKbV4sp0LEQwpOIQKRvBpedIE9CDlti2x6eLOupUAmKSZSdlHQaAJmMYzVpKNfFyKhFXgDU
1VKOQBvToqSqyMdYldRuWEOMzvqZ38olC7dVYfGh562RkV4gQRNR4DbdkvjKhpraJBwxlM9wzea0
Hav32BHvrvEezzh1ALo6JPYcQX7yEAWOZyzvUUNzRCAvaibB0OYBBfVsr0/564+67aGrAMymeZ8F
l+20AUYF4ifo8ZWygWuqtiIiJkJaLgrqQZwj+yBhzg9Mzdeto84VOCsSacJwE12El/8abkrbuqkN
giTXzJmk/Ylo7kzOg0u6C6DJwUDVx35jr9rfUS93PBnq8dF9X0I2MLk4KyAtLKF3AwVdzlbbbdHu
RcGUZTqBDVa8aQzziI1oAf/HVB+uvhFjz33HMLO69Wk8bLiwqGPGk05DXdTABV7M7wvt7SkQ5qrH
vJLmBHbSQW/n+sHV3t02JnhFOsoQJdT+S2wln4h61RFkuEzgsIsMHEYXyF0TrBMQAc0lBlR21aki
yaBqIGyyUaKbSlCZKeGRFoVqJxaHOhiNYa6cufUSDGaHFERPWth5tChUPz7xjsyL5mSNPVINFweV
QrMi8FH1XZlMQ9CdOVHbWBY/AZHTuJOB3hXAmOKX8yP0m4ORJ2HEVUZ/hn/74Mb5862N6hOzztRK
yqjVK4T2Nz7HgkyqWcdEl941ws5lvbshscO9yy6DJut7vDmXBwPdzHCyVXnYialG1xNy1LNjb0Y1
eVw+pQDkfAcmFvYUfExz2aD7K7PUwZdfZbgXIKSpNbfvmrn0YQd3hXbB0aqXRQ88D2tfyvPLdywf
sGfHyyZKCpJc/83GVRShwrXdE2O0L7KudOCbU+MCS7DMtNRtaCwd2snfVl6ljIfX//4hJqlrEk8P
EP2MwUWubG76GhNxIoJIK/uMlSRLzcD8E9a41go6H781UTsGGPnokNHyMhpxyJ4LPTrJWquOxJWK
MqMnLHrE4fQ4RdYFvHBXCrQdV9cB8ZBwwfmrk5yGwsNPtkSVHRX0Y7ECzIXLGR988fDKSLirDMNj
+3G+preZEDOv3lz0ALAqvVphrRPOvVaoyFhC7paAXzrbyt6g6tfrU620YtzafyQgqL7ovixYp2W0
xVHGz3mSS8qASpif1AsnzUweRv7eq8cuD2ZY2CMH+58Sog5eU3Opa4lvxTtdC40b1yuqgHSnTxHb
1P1SWbT9OPRNUxsqesV0eeUExj97qthy/y7SNUvAwL99mpsU34crdBOhuP2A8LZF6va872nmx08d
yuvG/30PFiAWfNrYtRc43Ur6FTC1JXMhCtpX6NtojIMIyDnccvEzY8P9HBQ5trmEHyvYEZjSMfbA
1p7DgV6bRuOJa1YEEcIRZrdsU6jgex7Bt5StjCVZE60ENKF3OM9UbznbMmd1FV7TqxTpmg+jRc/U
Ss5wY+LquieoVa6HhH2T4wm5e1ApzVa3k3RCi+6Cx0SnPav2PZ7f5Klk4JOOhMZUeQ6naa5ZdeZY
hG9GDEhWsi215uI1kbIKA3NBvS/K7d+KxMtM8UqU4XoxmHJ8G+6CXvj3p7NRyuly7WU5SIAfwqse
G1bZ4C6/aS7rLp9izZQJLsgQuumDcusSZLVrqLr8uNPQmWm5k8QpmQrs2N7vnEeBVmk15mQLij39
33Na/ZfyS7CrxuqzE3G8O+9vY0dvIlAv/Rp4cZpEeGcXQUEaYDuqbhpD9vQcN6HXuLhXhiz4BfHq
/ZuvvR8qPbl4XSq0DNJmPlaPHWqK8YTf+AgT7qP7pMtWhIGKtDHyAK8EAbT+OCtdBXZTZxXzZ70b
NHjFlyveoZ2FVeg7NTGzp+yaDSdu9di16aLQ1zToQC4VS/gHsY7IIxvUCSKkRPl61vHIkVKzMUmY
YDdow5pmXAe+zo+y95JDte26kEwtD0wgwxvAW5yArcblp4/MCu1YLvli6bX3yDdixqUHOA3Rw32B
BC2Kl5cOXofPhauzF1PUM5oe+r45AvW/ebf1ln5MMoBWkuYLqrZVZnet2zoxhpmlXDkFyaVtyb4W
WJ5nSF9+qva2soo14h5b8CEWOEi4CWvzlETJ+t2Jwc8FJ1Bqd6yj3oXPB1iamyOFosCRrkGC6Ziv
6ecXuEdEsfsi2HDcek4YwKHmY+kFp/g7b3oyRcjnOVfYDjDbkCBrm5zMEwuwrbSPbM1watmFhM8U
dKPmF2w4Q8NvP6cL2t1PkTFjKeOlp1iV2s6UmLKoj4c9SnyZThgNQki4JN0BxmsL8t4FUIKQP/7l
bTBJ6kt4LplL0pJzZrMpmk2Rav4rjsCBQQQkRGsFhmwQnMYuHcOKwUHoJOh+pMu6PIfHrS/m6EpO
YTovTDVir1AzqiIayb2b9EfG/iMTu03Hr37RiJpt0kMZzXMTDWV3TaanNftoxGFegckFM1m+V3hV
1tuFulVUlzSgDWDaFpGXdsvPTHyBYjJCAbsUMC5X7eG2fQ7epGKQ+Ye96E6b695hm6Hat5oJONrw
2Ln+SwgJlwDjeAcbLTbwiSOLQ+B0NuxlA3LcP3gP1xZLAlUPYtX4zWHBIwb9iHBYLVUhoxC2lkEJ
K6KxQmsJwrrKcNk0MF5noUIC76vD/4vH8BakpwQ8E2rPjCbO2pzIsj5Qj2qH1rTypfhZs+SpYRKS
QensWuf8PZx54pAkacmxioURiH4xr8X2TdDvdnamlQ36DZZcOuqLU2aX9h3H3OLOGe8L07EBvg19
X6u1hfVT3/F7guUObYCNWl83XlLLqNOE23BQFyrrNHAKQpEaHX/XlzU4q5XGhHYCGgW3PAauG4Tl
kBrJ24yadFHU1L5ByYCbzwZkubzpk8FvZvD4mq7qQq9ATiVn9jGsSKFtZx3XAS979V/58ozNQZoM
IzQkEvbMg21M7BtYfv0mQEgpZl0Opp0Z1TvPbkXYjJJ75VWg0BbLQahH/QWQJ1VkymW9IvmwSiGK
7WmXAvlwvFDzbCz2Q7sFmaMaAHHPpGYyXUgPAhQzOzuR5zHwbnV9MUDyUgQ56vkydKZjptWL3c+U
THqPgLVM52hpoZp24mnsw2Z8WiaeQtx/IU1G4zY0ZimYFFgKmHm2Ev0geg21nSS0LAwAcch5VC9S
/IJF75/o2c67WA/Cld8i1a0SG40j+4y9QklEIBYT1fg7MDp4sNnsAQE33bvhO8TPS6hgRmxfo+CL
6A4Y3MCVg+Hn1PNaWdwpKOEeSxy9fyZpTO0zy1XfZ/BUepnDsICoCdxlzn/0GLe6YjvTTjlvtwMI
uqZOLtJlN+gV4bPR95/+ij7mUsJh6HX7wzt+KRESSF5DNgchlxho4PR816VVys3cRK0FvNdANvr+
+dA6WknIdLunaOki51CRdsWvMNGDUwVr0CLF7Hx+SLXdIJuwgxM9p2xJbgrkuCI+g+sp6bb7c6G3
akcF0P9hatf5vpMhSRg4n/Lvf5nLMIInd/TeEtrCssqfZR9mOvBoeXdLxT7TIo49mBP4dqjVm6Bg
CQ7d/hjtIcsM2xnAtBrsZE5RQS02HZV/4zw3wsqX4SX6GTmlD9MYNVscvIGxBf91uh1ftKud3LgD
oL/x/lZkiblhsHiEDni7Bvcp5I8foBPMxa1RMlHRFE3t+7hp9s9GVKL+Mr6wjf3+e4oTGVnq97LE
VTiUKCxAVNSYahmcO208vUvJmE0VqMmor6lto+9WhRgTj1dvpbNTnxIykaF3ykpGpLHwXSYKb+6O
mAUNtzNT7Hhk+94YpY7WoX2/SyMREgwITqfqFsRwWrlLc7CnbYO5TT4A78QRpcvA2dri7xXyN58+
oYZ1041TUk1WUsLQ4mkg7Lv18sA1FS0E0vYjfNdA+NhCz7ReDEGrPYvJRUus3//vyrX2r7gVXaQE
ECWDJDwqaEUhOTS+19CWetz8U079r5PBlktSFdfI48ObDk4bVxvsRsMY4AbMiB1brhyFECMebC0q
kwZ3QiGShda6yc//3uAGpg8fFx0dI3j+/Yh6E0l074Y0HerO/vayLMz2EWv47DoJbTbz9IH4ilDp
K2uObjyz4/YaPgtF06rlsMtHQKDPOqcwVWKMoHXzvH//iSgPm5jIU+fI+3TCmK7fv9h6RVsIfG2D
zHS0uS0gmZhZgJ1PoilNogaYeuH/Y9It0xJGEiG+BgU355pleTn4FesTdHsl5pk1q2ktE0J1fi1V
TGkjY6k1nWc+riXJHBirWcUn2rSiB6BEbjfjxks+ZQmmgvjjiXxb1PpN9V1Vv/QJXEvDX/1dax80
Rf8OSz/bu2hUC8GWUl8f2kihgiVNFQQcOMLQhVfWfOq1lqO0pJRv/Yk+yTquSlo9d+sPfWthgKj0
Xf0EXQsyKhLcw7m8G+gjrNrniwDHthrZ0P3NkggEaSvASB2QgPeEkjj7W/x6eSMNcsCIYqHAjnQC
BxQqI4cyC+jjQzgDxRYd/5ejJHPDCc17RZtF23qFJ1ZC/hImoa2TmSNYvGbyNd7Ivsb5QLMiRnoQ
0NWb5/Bm2H324UV4Eatgh1DH4s7Dv9h3e0X6IWnB+tGy18PqzMbM1N3nvAUSQt2M3NJzP8wGLJS4
TJn4ptUnM3qq7B7hAW9HSAfijM0gvXovs/zDJjauYwPwjEtJNcHK8+yoOWCaTF0VyE5KMOV9mjRp
z5xKdB6nqRgZSHeZawiAwmbqZVTxBhHbOHFRqE6fIkjTNTrXkF7M7ZQMmtV8WkTP1AVunGYTya9b
x8g/llTX4HM0m+/ISks2CE32lRnAa61euEenB4Vn5R+AsAsxirFYaX5qBowJ9cY6vUR+8oK2xtNM
IOSqZroJmXupGq5r4qqkFuZCPgiIhyZKoM0Zk+Y10h0ax7w06fXcc+F0uhS2AtFLg2x/Zd6ulIjP
hwIuAA/OtGxZsoD2DKaUV/3P4HSrQG2GLMS3jAThAShihqmSX1fhvGOuyKcb99vRLY2h0+daHwas
JobCdqCWc1LbmuzIbB352Zi1D1rFo9k05deMk8+C23xEAvjp6gKOm3XN4boGdMCe0BKVZLNFS7nG
UEVyJ4H3gKPZSnKh59wu+Z+a+CAtWMoEIUe/g9kh7Ng54OS09wzJFVYSvpaNMOYPPV1vgQ2Y5oU+
sBNPcJf/+qbjNXJsOQbJl3Ep2QwE7VWLmtwAq8/cGH7CSg9wvOlmCciAb4ZjX3MDscWINqN/+sG9
F2m32c1ycnu2wi+0cC2MiQewTeaQ6WZozQmKvx67KgCKc/vGXJbyRF6pC6kNI9+PrGMImdQqsWAv
KmGh89mZIakORDK8mDGrtvV6/D9seNdf6SFS55Ync45OsnKZW8LtX9FqvrjnAGtsAgnI4XpkODc5
ODGyDAIk5NAPiK2ELWrM4l345QOD/UhA9pF1xmvUMVX83n4TJ9iyibOdLSYopv+bk2ymMk48BDbq
fNfPjtLHERFc3VAKTViVfhIPmcML52O9/SYA0Cj1EskEF14AtSDS7nqeyCwuFBJR9O0W6DdzWGMI
RRBJ1on9hI+iwUmx/CtgvppCVnIW/lc+4dey5atCtBntYvWtaHQPb0FLWU9pXmPPJlsRA/cRgRIC
7SExL/H1aH+gLf3Oh0eHUCBUpTkvVNbvsYL+69niDJC+RlA1VlHMf2p6vB1ckMFrWci34ybXkdBj
Ocr8zOzqVg/U0re2kQvdPZhV+jPwtMLWZg9PKgYIU40FMUtThSWzlEwYb+UMgxa9saKErWfTHL70
SSTnZjGBWTTMx2xnY89J71adXcmBbC6iQWUOqpCd5cqzQ2BKwFoX0JIZye+G+v3tY5KcSjsZ3XKT
snQwwU2Ja+cpWrkalulz5R6mPf5icHIvUl0KldAQ+LdEhQ4OD9FceoN3jn4vdO+/dZUpOqGE4vqm
F5cjqKLfbvFdaV/k9BpvBMAhgelGxq0mlgADOBEGFrlFBORFlIt+G5nCecl2zVAULTNwgnLDssfb
Kgb/Gqcj2tvXWilCm8zA0Zs7ct+i1E+XW3gT8GVOR7DOahC0d+yoD82gOsWIJ2DxL7Xgc7SZHQu1
PeuZ+Jcn89QdJfEyIDo0+wN3pMIinqlvuGeGplJjOmhHPj3EUcGdnyrALv0f2bE97KizNZkFK/U8
UcpLNQtSXd4uyVh+V1+OVv/3nvQsq1WFsc2VkiK8v6fX3cmn9DFlZB5UHKlz2yIQwrY9K4CwCSh1
bibSEJPmr1WBo/zz75+5srnJ52R/w17KL8wyq/n9hAnYgvHM5/OOUwpUhdphWKORtswmEH4AtpS1
3xdIu5dfYgzRK1gKak0/vx7aEquubNdR1wI1v6jONvoFJa3+8f/+UJ2WROGrn+buhBg+Ab9DJfsI
zu8yE0orMWdbCXEjRO3JR7Mjv+r1hC4mLMpM/j8DYMTpRQaNN02oKXaocu5618rWORke5xCbq0G6
YWWZJApe1Ssu3RN+9vCslR6esVTllgBa3uZEBE8QYXdI5naVlmmXJqT/rC1zNum1HLkkw1oRxO2C
bEvlhn9wTCJUPXbONDHa5VDS1Okd84Ai1KVg7BrA/BbJp6beWi+v1REeGzzybS8un37/6icmUhda
w+TVJtCHLo15VCGW00UPC2SjtPeBd1ZH8Ro5KPRe6c0Ke/i3urnqAk3Fin8lqQ+jJTp7PUVLzgNu
RRK6zIu4IqQ+qHckZbwvB3jVHZCtEqzqM74W9wJao8IP14BsxuGB4LAahdM2c2PISzVfgiA1W7AF
YlvgREwnYYhTOp/ilPCZkvodsLo9xAzk+9WGCYTjeEDKfO5vyo1GUKswJyj9Jdt71+qoTayjGzXb
AyDiZe+No22z4aTt4W3SuDxErAF6W5mP5g+yZ7W+Emv+JIyzDsb7WIuV2cAhhJ9q3iOAlzXXfFa1
5y27hzGFsmu85FMRVHhgX0Fdam3eajSSFqJAdnomoIQ95UYLTFlj9U3FuKUaFhFZuQrKvm8jcLYM
Vnxy+yW/X0rg5ylgQzaBgDcOzmzL6svbY9NiIOwFCbV4isAo2lGYH2+udlPGlyXSqw52ogVg7H/I
Aj1s+Nx/zycfUhtU+y0khh6Uw87iDPOuTWgT62vyXya5Ss/LCFjYZa3fTPrP2vkkZOSzRtEOI9l4
T0cU5aM608WFppMh4KbgIjqTeOp6B2/siiM6i6fVXUsnR9zIloHk0k8riZtOSvrW2H3xv/PzRNpE
RYCTMuPBQhF/zTvtzz/VLzLTWT+u+nIuFZypzwZj3kXP8+b1RfLVpEoccdJhCOR3W83gg4NRe/Dr
eIArmked8MEHqEMg1hriZCdTl1otjT8Gl1V8WxSmyUeHm0c8cSN+3HRPNKE5wNTdHPmL9bTvCVfL
VYkcfMksEKYII6WrgPW0SSXaIGpil/jsayAbnhyJp/3ms4Aw1XmuAFfImgyJ6cmAEqoVrA1Nx7/F
Z0lZepQEkxieQRRn3PP1c/3H54yDv2/FbjRu77hMO9jc29ZcKqjkp+bPuKZi/nHUWxH2XiLK2AQO
q/ai61eNMPfgVgHgjALEHMPq6O1AslbAMuixLS3Jxy8E9hvcqQSm+nt/h4/+wDf5pA0FjHaT/fu2
82dhsTRAJWLzPr/8UPsrLX25qPozC0lN7bjPl6QfHg9422g8eRGlk23/f/JzAyAc4iVBXnexeG8B
8mh0pGjRehTLcY3MmXcGCFxDfh7kfwl5ONlGKFxz9h57EKvN0uJn53qcpICqKxOT9C99tlb9BnAg
UTUyZjcpfcAChFK2M/bf9cqdX9SXsG4/PTid6OfTr2pQlCb5OPx+qey16w1ivC/MbTxxGELaS6em
k+y60dY5PKUa52J30Zb/jZrGhL5KilTr+6s0Tpvd4JqOX2TLHrH0rX07L+3/9cP35et+fcWTqLWu
8HJ/+EgktDrt9+oCzZpgVLTcVMoqPKT8sfZLwZPNuibFXSUqVG0y+/1uw7Ah9Ws9UJJmfNl33C59
UrShjuXiRLtxeuC8Y0PEz1FGw+1hBt0l4E52ama+dykivFPASS06oxgK2IL5MnEkvm7mJ9EC+SiH
q9IHeIrtXin1QqhfmLWJq2w1E39bak74nmVtrrvZEtgPpPawt3LjoBLMZ8lFtHs8lsxgLDGbHAUp
UfKsQ0XVKv29G5QWcUTUziykcouymxWTUqiUaIE6KCol1WlUQchhbQF3Fj54tZVQB+I8uhzNGnlu
Pr8Y773BJqv8onk5k8ZD9m/6vAcgsZIQj17hpgQAs3W1ItENoRZOEXW3X4uEHHejiWjPsSYtpHtg
rfLqhc/07PRaadUuZr4uhJGgXL/Mkbt8UOHc0AzZbDcF8MQ0uvpOqPoFE8iPpYpb+00/WrtJ6OQz
u5jaWC6dJkvdxOwR4auWUCQY+LerYPM8ZD5EVXVVwCDQ5wAsyWdU1gTExO2rryFqXLo72k7Iern1
CsaFl5dNywSuWKMMm+WtZnAevyYwb0qcQyU6gjPUCGH6ncbM2U9oYO02s8yBONXhBan0unqGVZlE
Zr9UrWd7R0p93AnXG4aR0YLnwrRHDKYp1HPwL7zrEx8ts5DVORXscM9Y16D/oDyesm/lqmQzI1uM
tdXDzJj7/VYUhk9cPieyQmn7MW0z6GBfY0oxDFXy/FOMhaBUs++cQzNFAzODx7iat974k2Auykxr
U9MmrRKN0VQzWOrXLLk9AEDqzOEezpsPEBtkxV+/ySY/pxEHXgO3FCGDcb82EYq4Sx0xAdvTtA13
0CObxOmdC0T8jUHOIo3RXQF9FMD+wMzeJ6EXbvrSEqBdfrmVq1ox/bZl4JQX6JeUB08xVg5k39lE
x+Ecggydlj+KMGtvH9CJnm8MX+zVk4t6On3y5/LpNKlfU7tYxLQpENe+0fr2Mbpykw/5Pc2FlDNU
qkhS6pryXk6hDbz5FY8LBUp+np2V+r6DbBpB6DCsoCZq+fBpX8gMgwLkffxuwYC2QtqyNUuoM9Rc
2XSlsfkwIKphY6cRGThauPiZ45X8ZIzbmpKtyWBrf1k42qYLs7diCzgNIipZq+B97/2Pwu3TKhHP
PKYP233zCcSzSHgTHUDkI3SBHiOeNjvYn8EGDz3A/xmGBK8XFiSDfYC6VpTfgycD/a5WWqJH2eUN
eRDMmaDny/S4NSq0rr3RYUKySRnCkDaHutXRmqq+2rEWKWiTRiForRxHBK4psGnQRJKwg3OOXUKn
qfLxBTQeOrdM2Na6cCQW/N0ycMMQZPE3Etij1t00F/qfz2vLfYsq+75KxZqr4avFJTG8QY5TnvgC
IpzOQLKlMOiq9rfQgqgOZIHTsF9PFEBWzAzC0Y3HhuE3ptxRIQuBcGRyis2kMqcBh1fPLVy5qb/G
QYeVG374sHX745xf4wqTnqtWoyHlIBOVr0pAEqfJQ7bj02XSZ/PTexxSXyTXa0d8GFo930tLZtMZ
bnyd7bNdioR6AMHBb+bvaoZI+wl0d/qvgrBQ2IdbnjnQoMZ6ML68AtRPlE+tVIEQ6ZVVgdunb1Fo
lcpihe3emml7JxRhFCMYqq/dL0kO8F6k0ok8yuu135FGITEHFNIXgrbBgPclcUbMUKQjzrwvCjjK
j67YsqweKmLc3hO86AG4mbiBw3Hgntb1J7uVvsQw0JznzMLQ9zUTcpoRKITGPkgns6pYonIkjv0V
5O8lCpqIT+0OKtxyLFAho2gXWqn6qnAJOWd1FWCTWCTrDnROU71KTTbaPa6IXU/owSP7wwzAkRxJ
f3ArRWe0fDAUhqcoJrFPMIbRuUNsPwYqgLW/zZ5hN3bVbbX1FcraC7vvQl+afOEfVxvi27YeycxK
WYnNLDlEiuP0MvqWi8FcxefBGVLWHn+sWfTJdt2OVmTKiizZzdRvV8BpCFiNwskSg+VPkvzQjBW8
b2i2DuLWr+kpy2p1eEAux0oxY/fYcO3U2vqWkjL01+fdNs3s2lndmBsNIeQRw80xZNrN2rk2zDFI
MqYDJPktgN7RKdao9Ff/YadJmxkjpZJ8Uoa4Q6PwGJIwnO5N6kEgVPv88lnkK0+KWKyOJL1LAu7g
OKYKvGbY09iDsefjSIGdY7A/pVHKHmOSHA/pAbcCT27fMK9Xq0NqfNx6VZd3SNiOqNiaHpM6u90W
VMHxHnZtY7R+PjdPsHIkk1vc+AQq2zY9izPEMehDqxa9jyIViKrr00arsGFLcBkJn6DXVKVbAHp/
JsWJX9Dea2eOp61oyk14CTlCU1iDoLtj582cJxClOuXADesRLRTAEwJykvQ1TjgV18GfmjncAJ0G
QrEv2QPoGemZz6+tHisM54D8EPelJaf7wwyXvekJO0Q9zo/0AUOULsAco7TaBXQWh7iNqAc5HQOw
E4wjvLpav/biM1ujObgSdlLjD3ZF3r6yv13NpT2+3ewj0kAY81E8ueCupvDgh+sWN5V7hFbfUTl0
n1OhbWE6sB6QA6yhFdWxizVdiVXuJ2u+1EHrWDffvhrjf/fWalTsyqzWW/4NLzXyLNNe54oRNaU5
Rp/DhDzArKC8cilnBCnzYKKMbZm+xixZYsgh7PakMC3G0ezo/v2+4Sp4+1078b1g4AGd/XLDl/F1
KJyC+EXhS510UJFnHjfUtjyB/Emffal43rcUTDHwW7kzUaG1NOFLJkA+t/SOMZCnPKlqnj8/LkYY
wfF+yGNEbH3jTCnIaNXNABUcqH4IuVwIdzR01hv0CYngNpIAi6DgRGLsUSxxonvQVv/TXH4IVEsG
3eEiohRwgIUOmkAisHj7jcbySPQ9LY9YjRdwuqNAekxoxPkWwfV+NuovbX9zCembpz2JB2UNwx2w
rnBBdVtsG8IcG/bOsu6Ad2ztxR2yY/PqdIDYLnsm9hn34jAnfV3w6au69fXBUE5ZtOiJrWcO5fq7
mj8w6F26d7ptN1iaNVAgIKFh81bWVA7whd1IscqiuNgCs6wIAbdCrOaJuWT2lBoRScnUfuserzkL
lmzqLHasqgq7132sobXw1xYU5tibhXy2pCM5LjX1hONh8DeDTYeqISRubYcw0NuaE5pLjPQUjr+i
91LrAmHZnknZgQ0RQVbOphZxF5m8zQaG/Ig8koNSjJygIffdJuCirjiG5Wyr5eM+4Qo51A0Fpvpf
KE6EcdeLbqo11epS8xs65Kr+ZSRWqH4EujN02A3Y01qPjIjwVWHGP4KX2u/78d8EYz2kwtHu67NP
ZHEPUW8ZVhNNwkj8AvyHmnOqq0JCSpZXP8hERBFGxG8rcTdV1YvTaMQTFDiFIfuZO5p5G85a6lb5
qJ4fC6qQ61N56kntvUgs/cxWix6kW3ne+rbywWJuYXULpLpzYnBmACzeK5yYzUbB/6NMrgtbAnuX
oeTLaU07VkBs/W1V3R9GPxtGy3E93hFUeXB5bpkGoB0RrZItxhbbUYDBF7ZcCPYZckg4GEVB1HlT
afVRc6ae7Ug+Ewu84oogdu2rq1vQTwlrUmV5I5834CRCKEK+V79jkYTYhRAFnPQ/kG0QwJgNtjA5
f3GPOgxspdIgJ77Bn3nvPLHzOrE1KZ7U2eJQbnQvkwozrguKgEpUZ4SRpTtUIj0XhLkqteKz/ySq
5ioeChrfKhdL7cbZ5SlHl9z0qhgWIh6/VUzMkDfVs0a4JTVxVxGUHOHehMJchoZeywDWHup0SMKF
jBar4tKlWLEnD8Fckd3ikPn/6IgUzJuTm8LqTZC3pOp7VtyuA+w1578DQ/Oio3I2+SD1I7LOmdmp
HWVPmaqXpmTHmsUX0Tb1y0UYBKDU57e5QLj6w83GlobU7Y7picc2EONtOlT3WbgL24Mi5v7k7Wec
wHSnm/En6jz51Sj4dpEQdKAwAPkOodPJg9r0VWYsR2/sgeOyGtBiCO3RIgn0/gUpN+xx7zKA6f0K
0cSwm1ZSgKspg6O2MDt4vWYW+8d4bP+8qmieQuLpyDV8VJdKuzaEQvng5JmIigsL45AxhH3spDG0
ZB4Y1t4qy9dMoY00VlFpKJ0uz97eNYO6O7t/UT4E+l9jf0dLtE5PoUQr1TefijqMm4HFTrJvqJLM
lsR5sEEVQfMaDoC5oMOUvhgulKSgDcrGLNcpY2tFaSsFLDJR0M9e9DLXhldVGc6zk27CguA0COwO
8TdFiwNArL6hNkKWMdsyglUDGjQQvXmJSKyM6vBG4fboPd+IpOTV8jjMb25rvkwWujJBpQrI4qoi
3ZAeqMaQ9y105e9MZ8m9hr47uN0rgMaBjGXx0rWdszJ2fELYZS6nsdsl9C53UcWR74YAV1BCi/Kl
P9EP2dR3OirmNrLkJhO3cJvY/nHRedTJogPRKdTa0GMD55GBCEeyv6/Bk+F0hfUTPnNwb7dKAu9Y
LoRhx1i21ZF2uEXEvqT9nvRl25mqTcyqUGqlVyq5/e3oy+Q9EUqXwnVdA8boR5w7eg6dEfGMbb/c
qaSpAKe1pGvoorNOV+Vt1u3zjNweRmedvCpENT4v6IQ8pf2WZQFGNrhzED1UNAtBAPnNpVBKn32Z
97L1ZJ+X2ZmP4VDRSAP0fmq+/X4PQjS2B6rQ7PEmDRtE7Oodv4aqpt+QAAzIm6dKIbJd1etFZHXc
eBulFBUIQfy01TJrfDvlJytSLNJC8KuLYUCuIh17glj6UQbNVf74pxAKcI401itxSOG9AB0M+UmD
hGfn6EALTA7mwJC/rXXPyHRjLoIMOm+ePfl5u/4v6cnt2EBEZNTJG13ZM1JHZl090//dDovFJ/LU
RNZySlxW4Y1f5fqE8PurOoitEpNqRpvTjMz5uFGiLLW7plZDeHNykSX7rdlMJGm5rFBM8mlpUwL+
+bU/pNmBC616wP3LsiXCc5ohvBFmLSBu0YHgHrolL0HDE2cFFl5vdxhKqSa0yhNnZ08MhQoTUf2E
DZvkoGR72jyV0DahrTMDR5iirIsoQslETeqSqjZpisf0dHCdf3vIWiSZYVqnE6wuPcfmf22w+8qb
16tlvNNbmLFeNjPkolWgBEQxL8JOeKvGl7wHTDncm0wTR3eXuILOLHxAldbW0vtIsFpQajjs6X2f
Yo+qq48rnbkABZh8mMAeE7bQaIqMfRPvaKKjA+ECUNZh3JWBxz5MjhmzknKXLQgUCkjLzG4J7Y6a
6/SZDydDxKLPtUSmv0rqknT6LhytZVy4gqquO5W+xka9HHfS3LBBnb+RdToZVxOvjntjsSwp/ICN
I4/TpE6+ZATa/5pzXMUsWzfrVtcHSPz4VU+HTspE0Bos3/LT5s4iC/QSISzG6H+cK9HzaIkmg3jE
hxWTsFyY8FMrFDViV5f9ft8+vz98UbDV1n+0BGRgPQpLM02zmbT0V7SXMlmoB/22/vGyyE8mEskd
m3jGylcqoACG4onoBdymhLWc2YMOrpGrADL5qYozx4qSD2U6JZ6M6khg8kcUhCgOTshy+4E9Go4O
ufxr+7Xnz8k14e+TR4tvcvMVj7samuu7kaZRL3Y26feIJIEmvi2Aoyz4i4Q5Nx+/jL0+GGhbZe49
lT6GJV3FuutfMbm0TS3nJ6TL6Dsf/eXt+503nzxW/cEtmiZ6ERUnMoWKQy5SIuY2SkD+LrDkxHNq
n8s4JniP38phq2gel3iPOkZm7+z9/jP+g9HjZRmHynLKaclopJmG7Q5SxOem5rk4OgI+jn0P7YQU
YJ7p0oePQ7igLXKfQckvXGCSvpY1hTDYsoHiswQZOy/6BxstOJBgkQuog9mBQWPzHDkHBWqMbQYL
uRMbkL9fRj7bot994c9d32r3ukpiccjPH9XveuU66ohqiIKWN2L3GKiSv/ACY8TpezgBPd4HP1Jk
/vfZkNkJ43rYoIb7gr0O8K0Pu2VDQVLVYIl+3g3JkkplU1GFKvnPc0h1pFl/Ys8TpQa2Cr3CiUjo
7MPNcNjgYuucLOSXruLJKEgvUc7F8t4WK1d8UogbEfzGKEYL0brb+i+rC+Icdzw2GhJaiMiMFqFf
KWDO3XlA4QDDjd6H3j1elqVzbLJ96pYOJswFEcVVtTFqrQzvuZJktSOevQGR2JymcW3hRlmsiBs8
4/fzrGToB7IJeVyq/bcFW/EPDDmdw1GvTSItrgPxrbPIDRG+HZuECzuHkDQFvOFXbHapJKu+PL0J
2oIDWUYqd9Bsy6jZ4HmZy7CG4K+JwwmSJxDZLmXkuoQgH1HfG0gue23xJgGf3me4xKGAySBvtA75
A23n+Vf9LLuVQ7X9Be29l6aorDsfc7m6bOdfW+lSFzrH+ApNbx7Mpf0Q8/cYuzkWjGemVICfNYI4
WoBencrs22A3NcS6+Rba6DovXygvE+M4Q4Y0E5SD6IzvrxfCbIfkolKCSd5ZFebm14Rn88hGzBtr
OkSRtT+Ps21G2xf7Of+tXyY6w4qHfohmxP+r0d5wIZhb4vvsovH2RgyCiuJm6QkKLVEHaEcFWTDI
BMqaVJ3Ha9uDb/nwJlyvCqLUeRBYqF1+agl7kuZi/RTx5bnHhOsoyBaqds0/S19TkBmmZzDpVl4b
JXPpq/7mIZyIFmpQluaumI3KQNDYAzymGCV1lrUhGrpn1Dp55dU3XV6WA15riFT3VbP9fssCA3V7
i/Fb6GPwx7WB1Tj3qMDohPAQR43rdYeoDHN00guu8o8FeyJRA4bRz1ddbbnD05SDJJzmPn3H8F3o
/CIOu6CKZm0X+mhEKVH7JtLBqaP0UfvePyXAkWhi3KHO6O1f9Ji+mbKVBmSDB0BGNQ1rZ0xIYo8Y
jnkCcxzlHFAyR+bpRzkMtelWgLYWcQ5yueYK03CLbj+uMNaQ7OwuL6Yma4BZ+0HsC6b4R/1bCJCD
tVtLd2ohpn1sFy0GbdZNOILPmGDlgqZ1uwpM0CLQ2GC61WwcDjYp/vdVwpMe1pi824PqezBpGVmC
SRJ3EccuXGHEw7weGmXn3lJulY3omrfAHwv88ZZWUi+Syu7Av8lc9CDksPgvcY8AuNwC3g9+dc5F
Xd5yaOyEDGZVatWMqQptdSRq2x9vyjnDLK+YplAPYfmeidL9rpUbsIph5GNT1l7JDbydcY2SD0IS
rChK97X00atsFfG9WelX7XgnNqqqhwoC3yNtFFQI58Y97LpSStJ1AJPh1ZbyGjL5lIfFnRrm/4Lg
QUiHME9jfPBAFRf4M9tjWV0YIOrT6r2qbYvTxUeKyrUp9TCDSW1NJIwmoijA5iryS+3LTkIfCelj
eiRGNaKAtS5YVMafAcihoZ70SFZkoQyDL0MfXzNURVFyyqrZTGp+gXeO3InRLS/sAqU6iDbOuQKu
quUUvh+tL6ibh/+KRXTNViybFMbJgdeOVWM869d+Ft5vFWxoHC3OmpJ44VNxYphAIUM5gmHqGiyG
fZY1D2Ao+NY6usECH1tTEDU59kD6EmM+c/NpRJCVpBAmjAi5SypY2Swye8TfWhD6izXNes4QBt+5
G9tjU9vH30zo16/14Z8R+BIVV9SA4jnWd6oh17/meUP07iwPvLjf5eG8aKnOMfRVPpxhhw5uUvNU
jjvgsfnWF4t/fZniFKTTDEK7dpOC3A+z91X8EorPFr9yM3WmQC0tx/dSJi6y1aDeZpcpvm7BJ7It
y96BlCpnjz55QTK/vy6EYy4SaVp4LoxeACTVVWzo+8QDwtt7z/3I/il6DOFlWdzLNC3pyeqchAVz
1GSpmeFbkqENJGbv4kRn8H7puNdEf1Pkm88VozXMjcZ3fcP0GmwPjy70CEp9DlpF1Cpa8HQAPBeq
IA4rXmsZRUmbG/3i+hxnFf3jSCrVOoPCnt8D7a85ZOpTq+b25aKwqOQbCanqptUc2yfDmfd03J99
AM3jGeS7fy2oynTgPH4vu6gq91SPdccnp3sOauvSU0VE7CsVYSUG2WDjo7Bx1lYwERanyKMmVTJC
AQGeu2/Ge+CX2HOa1qTKjriqqV/Sr2WycLR+k4IQjF5ITIlbQTpPTnDoh1jmWq8Sfv1jKUTf+Y8g
l6ng/9AEfcJPTj3OAnx8CQYjMmImHuZfrUKvkWGY3r9iy8AsWcOyy3uMXVKxEdkPREBvhOx1TJBv
SdTJbpU+sJMWTtCBOAsuT+Ik1eq9kHPIuG6i2on9wEiSERToN0J4U6SDIUA2qu6q2hN06gGKNc8N
9kq2CkSG0eim0xwtdU7a+NKKd6pPeUTSWA4wh30s+uqdpmwwxlQ/TXedQw5lqtLGGzO2sjSumZ63
rT+DH9aAAWHbMCsVjdDJ8dijjcnd3uh/2OivyQ9WxNS6crqODhJ5rDZN0fCGZkFap4T/323bgRTh
csSJgHXjDCVGrXz1Sd4NOZe49pt0Uc2ChpJmQQVHOJqukzZgM/ujTkWUDvkNWsrukLWqK2QRm/0E
R3P0qoVRZPXnNhnSepkyRn+MP9wTSywoNR0IDCZDSYWixK/XKiOV7S5iSxndKL+D2aPiaxNvcsx9
68EMa9kB8dBTJfTpNN+oMOkMSu8soA+hbL6WffF+pFxGsEkTgQXIIHsqNi13OPV4HnSTA4X841Ml
1QwQvCDwvlwisBP1xL3jynLKeOwsMH4ORRQWCTztHsLXzchmc2ZMhWoDVv2udyW4hKauvujAXwd0
RSX+n6K+VXHUHXMEFPm8Hk4fQhZqKsQnldqKKTaKM/V/9R71L7CbvxUOqtKrQ+EFZr0FGxDtcitU
Hc161yybbDesXztCwNLDBmDHNkdKjROhMrGJ53BjsvuH/rL2GKfqmojAc1JmSrbsMPwhRd7GXxgi
Lj80OVxGkuCve0+zyNQi7VV0q2x/oVywUz3XS3Q8j2yb57xJudY1vf0I0jwOuvXNblYuXodOErcr
alljezsD89c1xabd4L+Kq9nvhoxvlBnk7aOQ0HphvP6QWWHwx0sOTLyXRrCnDFc1qVxqyAjKCPHX
kvtHHwgRj5XygPRJUEPl3hGmg0fyuJUaq0w1VQLbXSEMAGP7FIm9VeOkWCOjewr1/C2kXRtEyRKx
yr6isgH9f1kmTmr93+P6IsCzy/br/vnYDdS/nmFwyo40f91x31xadE+KpdqveHqM/vDkdbR9NoMq
tc5AXhfbPhlyIkE1WD7HGVoLBlHnwBfDY9ZmMO3rM3+qh4teA321zr+Ug3f6Jx6h3yUp+La7raP5
rmkCyTaw0vpTc5YILfCgIAqgnRSATk/ETBfk68Yf7kXz2FZEOnX9lQ0Uaa+uiaS8J+22aKGyZm98
rilqVpyzF+ZVdriyP+Ge7OQpqwKQazi0sOcZd5IXkmhw6scY/maI4wIw8ti7bi9wqDurwumyDMtK
xPO+pWiAjaa8ZiQQqc+mn+MDrkz1li0IO/p6UqSIw5iIpRL6m3ltXEmRoTBCnmv0j9zc0irK1x3H
tz9O0itApA1c0bhial8XRA7lrw9XE5MvGWxpsmvpx/Eqwc4m3RJpYll9xsMhypoKXaK4YAYjnptP
bcNifiEkRxxFfeiXjnPXzhxWA3Q8a75WPVFaXFzaG0APKm9V943FjKYkwPcuUSVqnAVwxNw0MHbJ
mZGhiyUz4LxKPdowidvbQE/fsgfszGKHxFNJlsNRXkUO1sDYCugRv1HOeTmnXU6xvbd5XA2Q+ELS
KbBZERuPZ2alMIShXG3B0RuWYm1P9EKmAmjL6xV5dnafjPbuMrZhpkkOIoPfBWcHCduXQwmoIla3
65N4/n/U8kGPUp6bKRvfp/efoFpL10NOPo+e/GWG6bQZ0Lk4rjo5S1a0+I2gPmuROXTtZlDMzLWM
dEzsGla/WbLayjzC4Jx9hZGTlmVYTiB5UhKPsw+OB0r+ufORxlDNtBlmShfVoOSYglN4n7ZIhoON
ieKRZd/07Kbo9gIsPlmpuwvcSCi0MjDGpWpMclLTBBpYLFaIQtWIk088SJ1y165dgQ5Bm+UfENvX
iurQWR95LthJQ2CvP65f+et84JHzrvSXdN6J817cFJ+2PKgx9xgpmy4wyQxzIb3ki386idqSsKIX
CKs14b5IbOltcDQGLQdC9PriASCm+JiC+MEmJ/vkrl55SwzaoWo/b9TiHotyNMWPzQdu994nwpqo
VVJeXtplrgLtI0Sgo3olvuFnXY+Uz5j5i++1Nd8OEgcbVP/+/pTBgKxSWR6M0/i36mlDcA5vG4M1
bMzj41yHZCGHRooU9FJwVVTxj7R+03y/bgLxkGor8Q6vhQ30w+Zghxm3c67OvJnRJFMi1+XUB+LJ
zLpHZpfFTX0sHq1hAIskdREeNe4HylFSn9dNwEZk2muIxJEq9fXMVNDTjPpbYRe8vYZdgbGiedA4
BvuODzAV4tev/dGOrAnIoORSOBHwk2VZJQeS/7vKh1D7rW0xFENFKTYgbuaT53NOmP82sODLlMC3
TW6wxOJVUgTWE8ZVXJ3nk0jLvVeAXSklSd6aQIOnRVL1TqRY03NbdqpACe6p1U/hinzn3pJTUbGG
J36Rmc0vmwSB4nbvRe2vcSXzLJA6WW5quFuv9xLwFr3A0YTuJeOH6jBzRe+xbN1Bk2PlvMd65sua
9yJt7Um0rbqp29rnpDAewE7GkB8btHQm/Grrr5usU7V/lQ7GSAnqF7uATJeIm7oomxQhIVXP6Bj0
Qb5Rz7DO6vZ1CJbrnW/YBw4o1dVB3mBqtWlqfXICB9fUCWyXXX7IYd5ea7eLK5jeDf+QBwxNrrWV
NYtw3ETGSTT7j0c6Jb0R8Xc46VSoFG1U5MK0GSbpHlJ0b1zVoa8fDCbe3nVtiPuyGdPx1cPQp0pT
0ccrchdQ14ckduw2IM9AtchefThzNo+nGiNtbazQ5HpT4+JDlg6aGugV9+AMZR43zqpemdtaXLi0
3pvoJjDYbnuAvr7kWrNXaOiXFlf49WPMyB9UTQ30bVa+ujbxPjR4ztUT9FIhzLs4dtpB6oGs0Dl6
3feM3nlbtOWWJ/s9lGyKwYer7Zu6R2RrTYkCAUtM5e8Gawevb9rrRl2lSyn+zDUa595EFRR4GoWu
dnwSfpIPST2WNI4aZsyinl04xQKdC+OZyTnN+1MXmN1j9eQ7tBci3LpQ3ibxMYcXD7Q4Fj/z0USQ
uPRKYPlW9GmOPb1mr+ncbIeLnh2O7QaR1/EmwU5OxbZKs/JtKaMenxqVz4ssS48MT4Xegtebl7N8
MEBih2WhZQwEgknOHxvxZxRDpP7ctaQOs64RtNwzm+cvkndAKpEDkDvPYcWHHxylLUqYepKQasl4
bE5UX8jCwzmOeU6N6ecXXkeu6Pv+HuSmXJHgNLGL9wnYOJdYxSSnXsJGKqPqkp67Wi0k6WwkpB4J
+y4Xeyest5vRWOD+LTpUt0s8fLsJDiX50bRPLIx5XZr8m2n/MIyePp0Koa3UWam2q//iW1SiQeVL
TDK/LizD9xqWl7B5L6BAGvqR6yg1DrNOE4byoV9dIYakvS3iDDcF4Acc6nFc10KzFkNwfv/iooPe
LpZsQh9GF/47+wLGlxUNKGazzEaGvq2cwNLxcQYPPUSJSvDynKcijVqYSbFjhD2lmLw9m2riDap+
cdIoeSb17tQOyDAbufgDuJxALJKpUk4SOXkaUYJV9c6lfkVO7sXpGM8rTSxsx29lqQrhM3G0kGcR
Ob4mDb4Gcy6KIlQBTpnInak34gC3FOkJUdmvRR79SBUp9/VzwnuNU9fi/4xbXfyAuE2CCqDv4ZAC
RhVaYqvDXKx0aarhPFH8iaEwPm3YNi+ARsXD1EjibpCF+hWucYBjWNqfGi7EzW64pDmH1P7aMFMB
mKWx1K17H6StZmaLYWBoh2DObqf9MngeYGJDTd4E4mQtFWS09tb+zzhF1aciauGPShOWEhbU3jDI
3Cd85uWEsIzlTJeNySY+XbRwdWPHt3y7h3d7m24yXhxgFUogrA/9wOJDuAUh0V5lOoofRMnnpZmP
uzExqH450E3ZWDhjpc5VBuSmshIC9qBbuud9UhJX1G3f7q8WZRam0M+k4U10EiQUgIrmvIpVkZI5
ZpZcBssDay+wpr4ZRjvi3XWxdym4JBZldTGgIFG3CYs2UiaxQss6g0kk80m3CNce
`pragma protect end_protected
